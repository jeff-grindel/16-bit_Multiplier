* SPICE NETLIST
***************************************

.SUBCKT INV in gnd! vdd! out
** N=4 EP=4 IP=0 FDC=2
M0 out in gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07 $X=210 $Y=-180 $D=1
M1 out in vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07 $X=210 $Y=800 $D=0
.ENDS
***************************************
.SUBCKT SP_AND3_DR !C !B !A out out_b gnd! vdd! C B A
** N=18 EP=10 IP=4 FDC=22
M0 15 C gnd! gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=5.3325e-14 PD=8.2e-07 PS=9.35e-07 $X=-1085 $Y=-715 $D=1
M1 16 B 15 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=3.78e-14 PD=8.2e-07 PS=8.2e-07 $X=-705 $Y=-715 $D=1
M2 4 A 16 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=4.1175e-14 AS=3.78e-14 PD=8.45e-07 PS=8.2e-07 $X=-325 $Y=-715 $D=1
M3 6 !A gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=900 $Y=-715 $D=1
M4 8 !B gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=2530 $Y=-715 $D=1
M5 14 !C gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=4030 $Y=-715 $D=1
M6 17 6 gnd! gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.835e-14 PD=8.2e-07 PS=7.5e-07 $X=5675 $Y=-935 $D=1
M7 18 8 17 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=3.78e-14 PD=8.2e-07 PS=8.2e-07 $X=6055 $Y=-935 $D=1
M8 out_b 14 18 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=3.105e-14 AS=3.78e-14 PD=7.7e-07 PS=8.2e-07 $X=6435 $Y=-935 $D=1
M9 4 A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=1.935e-14 PD=5.85e-07 PS=5.75e-07 $X=-705 $Y=3505 $D=0
M10 vdd! out 4 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=115 $Y=3505 $D=0
M11 6 !A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=900 $Y=3505 $D=0
M12 vdd! out_b 6 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=1720 $Y=3505 $D=0
M13 8 !B vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=2530 $Y=3505 $D=0
M14 vdd! out_b 8 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3305 $Y=3505 $D=0
M15 14 !C vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=4030 $Y=3505 $D=0
M16 vdd! out_b 14 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=4850 $Y=3505 $D=0
M17 out_b 6 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07 $X=5675 $Y=855 $D=0
M18 vdd! 8 out_b vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=6055 $Y=855 $D=0
M19 out_b 14 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=2.52e-14 PD=5.75e-07 PS=6.4e-07 $X=6435 $Y=855 $D=0
X20 4 gnd! vdd! out INV $T=6065 2910 0 0 $X=5615 $Y=2395
.ENDS
***************************************
.SUBCKT NAND2 A gnd! B OUT vdd!
** N=6 EP=5 IP=0 FDC=4
M0 6 A gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07 $X=210 $Y=-360 $D=1
M1 OUT B 6 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=2.52e-14 PD=5.75e-07 PS=6.4e-07 $X=590 $Y=-360 $D=1
M2 OUT A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07 $X=210 $Y=670 $D=0
M3 vdd! B OUT vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14 PD=5.7e-07 PS=6.4e-07 $X=590 $Y=670 $D=0
.ENDS
***************************************
.SUBCKT BE_Cell Yj+1_b Yj+1 Yj_b Yj Yj-1_b Yj-1 gnd! vdd! TWO_b ONE TWO ONE_b
** N=26 EP=12 IP=39 FDC=82
M0 26 10 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.025e-14 PD=6.4e-07 PS=5.85e-07 $X=37275 $Y=-5030 $D=1
M1 12 23 26 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=2.52e-14 PD=6.65e-07 PS=6.4e-07 $X=37655 $Y=-5030 $D=1
M2 13 Yj_b gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.025e-14 PD=6.4e-07 PS=5.85e-07 $X=37745 $Y=-13095 $D=1
M3 15 Yj-1 13 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=2.52e-14 PD=6.65e-07 PS=6.4e-07 $X=38125 $Y=-13095 $D=1
M4 17 11 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=38905 $Y=-5030 $D=1
M5 19 Yj-1_b 13 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=5.445e-14 PD=6.65e-07 PS=9.65e-07 $X=39755 $Y=-13095 $D=1
M6 24 9 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=40535 $Y=-5030 $D=1
M7 21 Yj gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.025e-14 PD=6.4e-07 PS=5.85e-07 $X=41025 $Y=-13095 $D=1
M8 22 Yj-1_b 21 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=2.52e-14 PD=6.65e-07 PS=6.4e-07 $X=41405 $Y=-13095 $D=1
M9 25 Yj-1 21 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=5.445e-14 PD=6.65e-07 PS=9.65e-07 $X=43035 $Y=-13095 $D=1
M10 12 23 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=37275 $Y=-1635 $D=0
M11 15 Yj-1 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=37745 $Y=-9700 $D=0
M12 vdd! TWO_b 12 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=38095 $Y=-1635 $D=0
M13 vdd! ONE 15 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=38565 $Y=-9700 $D=0
M14 17 11 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=38905 $Y=-1635 $D=0
M15 19 Yj-1_b vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=39375 $Y=-9700 $D=0
M16 vdd! TWO 17 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=39725 $Y=-1635 $D=0
M17 vdd! ONE_b 19 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=40195 $Y=-9700 $D=0
M18 24 9 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=40535 $Y=-1635 $D=0
M19 22 Yj-1_b vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=41025 $Y=-9700 $D=0
M20 vdd! TWO 24 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=41355 $Y=-1635 $D=0
M21 vdd! ONE 22 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=41845 $Y=-9700 $D=0
M22 25 Yj-1 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=42655 $Y=-9700 $D=0
M23 vdd! ONE_b 25 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=43475 $Y=-9700 $D=0
X24 12 gnd! vdd! TWO_b INV $T=42665 -2230 0 0 $X=42215 $Y=-2745
X25 Yj+1_b Yj Yj-1 9 10 gnd! vdd! Yj+1 Yj_b Yj-1_b SP_AND3_DR $T=25560 -12380 0 0 $X=23610 $Y=-13600
X26 Yj+1 Yj_b Yj-1_b 11 23 gnd! vdd! Yj+1_b Yj Yj-1 SP_AND3_DR $T=25560 -5140 0 0 $X=23610 $Y=-6360
X27 24 gnd! 17 TWO vdd! NAND2 $T=42855 -4890 0 0 $X=42405 $Y=-5535
X28 25 gnd! 19 ONE_b vdd! NAND2 $T=44890 -12955 0 0 $X=44440 $Y=-13600
X29 15 gnd! 22 ONE vdd! NAND2 $T=44890 -10165 0 0 $X=44440 $Y=-10810
.ENDS
***************************************
