* SPICE NETLIST
***************************************

.SUBCKT GREY_CELL !Gi-1 Gi-1 !Gi Gi !Pi Pi !G G gnd! vdd!
** N=16 EP=10 IP=0 FDC=18
M0 14 !Gi 7 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07 $X=1045 $Y=110 $D=1
M1 14 !Gi-1 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07 $X=1915 $Y=110 $D=1
M2 gnd! !Pi 14 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14 PD=5.7e-07 PS=6.4e-07 $X=2295 $Y=110 $D=1
M3 gnd! Gi 9 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3125 $Y=110 $D=1
M4 15 Gi-1 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.88e-14 AS=2.025e-14 PD=6.8e-07 PS=5.85e-07 $X=3935 $Y=110 $D=1
M5 11 Pi 15 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.385e-14 AS=2.88e-14 PD=6.25e-07 PS=6.8e-07 $X=4355 $Y=110 $D=1
M6 16 9 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07 $X=6395 $Y=2680 $D=1
M7 G 11 16 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=2.52e-14 PD=5.75e-07 PS=6.4e-07 $X=6775 $Y=2680 $D=1
M8 !G 7 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07 $X=6815 $Y=-60 $D=1
M9 7 !Gi vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=675 $Y=3505 $D=0
M10 vdd! !G 7 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=1495 $Y=3505 $D=0
M11 9 Gi vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=2305 $Y=3505 $D=0
M12 vdd! G 9 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3125 $Y=3505 $D=0
M13 11 Pi vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=3935 $Y=3505 $D=0
M14 vdd! G 11 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=4755 $Y=3505 $D=0
M15 G 9 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07 $X=6395 $Y=3710 $D=0
M16 vdd! 11 G vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14 PD=5.7e-07 PS=6.4e-07 $X=6775 $Y=3710 $D=0
M17 !G 7 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07 $X=6815 $Y=920 $D=0
.ENDS
***************************************
