** Generated for: hspiceD
** Generated on: Sep  4 19:52:56 2013
** Design library name: my
** Design cell name: MULT_TOP_v2_test
** Design view name: schematic
.GLOBAL vdd!


.TRAN 1e-9 200e-9 START=0.0 SWEEP DATA=D

.OP

.DATA D
+	X0_	X1_	X2_	X3_	X4_	X5_	X6_	X7_	X8_	X9_	X10_	X11_	X12_	X13_	X14_	X15_	Y0_	Y1_	Y2_	Y3_	Y4_	Y5_	Y6_	Y7_	Y8_	Y9_	Y10_	Y11_	Y12_	Y13_	Y14_	Y15_	!X0_	!X1_	!X2_	!X3_	!X4_	!X5_	!X6_	!X7_	!X8_	!X9_	!X10_	!X11_	!X12_	!X13_	!X14_	!X15_	!Y0_	!Y1_	!Y2_	!Y3_	!Y4_	!Y5_	!Y6_	!Y7_	!Y8_	!Y9_	!Y10_	!Y11_	!Y12_	!Y13_	!Y14_	!Y15_
**Delay Testing/Verification Testing/Dynamic Power Testing
**+	1.1	0	0	0	1.1	0	0	0	0	0	0	1.1	0	0	0	1.1	1.1	0	0	0	1.1	1.1	1.1	1.1	1.1	0	1.1	0	0	1.1	1.1	1.1	0	1.1	1.1	1.1	0	1.1	1.1	1.1	1.1	1.1	1.1	0	1.1	1.1	1.1	0	0	1.1	1.1	1.1	0	0	0	0	0	1.1	0	1.1	1.1	0	0	0
**+	0	0	1.1	1.1	1.1	0	1.1	1.1	1.1	0	1.1	0	0	1.1	0	1.1	1.1	1.1	1.1	1.1	0	1.1	0	1.1	1.1	0	0	0	0	1.1	0	0	1.1	1.1	0	0	0	1.1	0	0	0	1.1	0	1.1	1.1	0	1.1	0	0	0	0	0	1.1	0	1.1	0	0	1.1	1.1	1.1	1.1	0	1.1	1.1
**+	1.1	1.1	0	0	1.1	0	0	1.1	0	1.1	1.1	0	1.1	0	0	0	1.1	1.1	0	1.1	0	1.1	0	1.1	1.1	1.1	0	1.1	0	1.1	1.1	0	0	0	1.1	1.1	0	1.1	1.1	0	1.1	0	0	1.1	0	1.1	1.1	1.1	0	0	1.1	0	1.1	0	1.1	0	0	0	1.1	0	1.1	0	0	1.1
**+	1.1	0	0	0	0	0	0	1.1	0	0	0	0	1.1	0	0	1.1	0	1.1	0	1.1	0	1.1	0	0	1.1	0	1.1	1.1	0	1.1	1.1	1.1	0	1.1	1.1	1.1	1.1	1.1	1.1	0	1.1	1.1	1.1	1.1	0	1.1	1.1	0	1.1	0	1.1	0	1.1	0	1.1	1.1	0	1.1	0	0	1.1	0	0	0
+	0	1.1	0	1.1	0	0	1.1	1.1	1.1	0	1.1	0	1.1	0	1.1	0	0	0	0	1.1	1.1	1.1	1.1	0	0	0	0	0	0	1.1	0	1.1	1.1	0	1.1	0	1.1	1.1	0	0	0	1.1	0	1.1	0	1.1	0	1.1	1.1	1.1	1.1	0	0	0	0	1.1	1.1	1.1	1.1	1.1	1.1	0	1.1	0
+	0	1.1	0	1.1	0	0	1.1	0	0	1.1	1.1	0	1.1	0	1.1	0	1.1	0	1.1	1.1	0	0	1.1	0	0	1.1	0	0	1.1	1.1	0	0	1.1	0	1.1	0	1.1	1.1	0	1.1	1.1	0	0	1.1	0	1.1	0	1.1	0	1.1	0	0	1.1	1.1	0	1.1	1.1	0	1.1	1.1	0	0	1.1	1.1
+	0	0	0	0	0	1.1	0	0	0	0	1.1	1.1	1.1	0	1.1	0	1.1	1.1	0	0	0	1.1	1.1	1.1	0	1.1	1.1	1.1	0	1.1	0	1.1	1.1	1.1	1.1	1.1	1.1	0	1.1	1.1	1.1	1.1	0	0	0	1.1	0	1.1	0	0	1.1	1.1	1.1	0	0	0	1.1	0	0	0	1.1	0	1.1	0
+	1.1	0	1.1	0	1.1	1.1	1.1	0	0	0	1.1	0	0	0	0	1.1	0	1.1	1.1	1.1	0	0	0	1.1	1.1	1.1	1.1	0	0	0	0	0	0	1.1	0	1.1	0	0	0	1.1	1.1	1.1	0	1.1	1.1	1.1	1.1	0	1.1	0	0	0	1.1	1.1	1.1	0	0	0	0	1.1	1.1	1.1	1.1	1.1
+	0	1.1	1.1	1.1	1.1	1.1	1.1	1.1	0	0	1.1	1.1	1.1	0	0	0	1.1	0	0	1.1	0	0	0	1.1	1.1	1.1	0	1.1	0	0	0	0	1.1	0	0	0	0	0	0	0	1.1	1.1	0	0	0	1.1	1.1	1.1	0	1.1	1.1	0	1.1	1.1	1.1	0	0	0	1.1	0	1.1	1.1	1.1	1.1
+	0	0	1.1	1.1	0	0	1.1	0	0	0	0	0	1.1	1.1	0	0	1.1	1.1	0	1.1	1.1	0	0	0	1.1	1.1	0	1.1	1.1	0	1.1	0	1.1	1.1	0	0	1.1	1.1	0	1.1	1.1	1.1	1.1	1.1	0	0	1.1	1.1	0	0	1.1	0	0	1.1	1.1	1.1	0	0	1.1	0	0	1.1	0	1.1

.ENDDATA

.MEASURE et_s0  TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s0) VAL = '0.55' RISE = 1
.MEASURE et_s1  TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s1) VAL = '0.55' RISE = 1
.MEASURE et_s2  TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s2) VAL = '0.55' RISE = 1
.MEASURE et_s3  TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s3) VAL = '0.55' RISE = 1
.MEASURE et_s4  TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s4) VAL = '0.55' RISE = 1
.MEASURE et_s5  TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s5) VAL = '0.55' RISE = 1
.MEASURE et_s6	TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s6) VAL = '0.55' RISE = 1
.MEASURE et_s7  TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s7) VAL = '0.55' RISE = 1
.MEASURE et_s8  TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s8) VAL = '0.55' RISE = 1
.MEASURE et_s9  TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s9) VAL = '0.55' RISE = 1
.MEASURE et_s10 TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s10) VAL = '0.55' RISE = 1
.MEASURE et_s11 TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s11) VAL = '0.55' RISE = 1
.MEASURE et_s12 TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s12) VAL = '0.55' RISE = 1
.MEASURE et_s13 TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s13) VAL = '0.55' RISE = 1
.MEASURE et_s14 TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s14) VAL = '0.55' RISE = 1
.MEASURE et_s15 TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s15) VAL = '0.55' RISE = 1
.MEASURE et_s16 TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s16) VAL = '0.55' RISE = 1
.MEASURE et_s17 TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s17) VAL = '0.55' RISE = 1
.MEASURE et_s18 TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s18) VAL = '0.55' RISE = 1
.MEASURE et_s19 TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s19) VAL = '0.55' RISE = 1
.MEASURE et_s20 TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s20) VAL = '0.55' RISE = 1
.MEASURE et_s21 TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s21) VAL = '0.55' RISE = 1
.MEASURE et_s22 TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s22) VAL = '0.55' RISE = 1
.MEASURE et_s23 TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s23) VAL = '0.55' RISE = 1
.MEASURE et_s24 TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s24) VAL = '0.55' RISE = 1
.MEASURE et_s25 TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s25) VAL = '0.55' RISE = 1
.MEASURE et_s26 TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s26) VAL = '0.55' RISE = 1
.MEASURE et_s27 TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s27) VAL = '0.55' RISE = 1
.MEASURE et_s28 TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s28) VAL = '0.55' RISE = 1
.MEASURE et_s29 TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s29) VAL = '0.55' RISE = 1
.MEASURE et_s30 TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s30) VAL = '0.55' RISE = 1
.MEASURE et_s31 TRIG V(PC) VAL = '0.55' RISE = 1 TARG V(s31) VAL = '0.55' RISE = 1

.MEASURE pc_s0  TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s0) VAL = '0.55' FALL = 1
.MEASURE pc_s1  TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s1) VAL = '0.55' FALL = 1
.MEASURE pc_s2  TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s2) VAL = '0.55' FALL = 1
.MEASURE pc_s3  TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s3) VAL = '0.55' FALL = 1
.MEASURE pc_s4  TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s4) VAL = '0.55' FALL = 1
.MEASURE pc_s5  TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s5) VAL = '0.55' FALL = 1
.MEASURE pc_s6	TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s6) VAL = '0.55' FALL = 1
.MEASURE pc_s7  TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s7) VAL = '0.55' FALL = 1
.MEASURE pc_s8  TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s8) VAL = '0.55' FALL = 1
.MEASURE pc_s9  TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s9) VAL = '0.55' FALL = 1
.MEASURE pc_s10 TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s10) VAL = '0.55' FALL = 1
.MEASURE pc_s11 TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s11) VAL = '0.55' FALL = 1
.MEASURE pc_s12 TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s12) VAL = '0.55' FALL = 1
.MEASURE pc_s13 TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s13) VAL = '0.55' FALL = 1
.MEASURE pc_s14 TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s14) VAL = '0.55' FALL = 1
.MEASURE pc_s15 TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s15) VAL = '0.55' FALL = 1
.MEASURE pc_s16 TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s16) VAL = '0.55' FALL = 1
.MEASURE pc_s17 TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s17) VAL = '0.55' FALL = 1
.MEASURE pc_s18 TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s18) VAL = '0.55' FALL = 1
.MEASURE pc_s19 TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s19) VAL = '0.55' FALL = 1
.MEASURE pc_s20 TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s20) VAL = '0.55' FALL = 1
.MEASURE pc_s21 TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s21) VAL = '0.55' FALL = 1
.MEASURE pc_s22 TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s22) VAL = '0.55' FALL = 1
.MEASURE pc_s23 TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s23) VAL = '0.55' FALL = 1
.MEASURE pc_s24 TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s24) VAL = '0.55' FALL = 1
.MEASURE pc_s25 TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s25) VAL = '0.55' FALL = 1
.MEASURE pc_s26 TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s26) VAL = '0.55' FALL = 1
.MEASURE pc_s27 TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s27) VAL = '0.55' FALL = 1
.MEASURE pc_s28 TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s28) VAL = '0.55' FALL = 1
.MEASURE pc_s29 TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s29) VAL = '0.55' FALL = 1
.MEASURE pc_s30 TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s30) VAL = '0.55' FALL = 1
.MEASURE pc_s31 TRIG V(PC) VAL = '0.55' FALL = 1 TARG V(s31) VAL = '0.55' FALL = 1


.MEASURE TRAN avgpwr AVG POWER FROM 0 to 200e-9

.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
+    POST

.INCLUDE "/home/jgrindel/apps/FreePDK45/ncsu_basekit/models/hspice/hspice_nom.include"
**.INCLUDE "/apps/FreePDK45/ncsu_basekit/models/hspice/hspice_nom.include"


** Library name: my
** Cell name: INV
** View name: schematic
.subckt INV in out
m0 out in vdd! vdd! PMOS_VTL L=50e-9 W=180e-9 AD=18.9e-15 AS=18.9e-15 PD=390e-9 PS=390e-9 M=1
m1 out in 0 0 NMOS_VTL L=50e-9 W=90e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends INV
** End of subcircuit definition.

** Library name: my
** Cell name: NAND2
** View name: schematic
.subckt NAND2 a b out
m1 net16 b 0 0 NMOS_VTL L=50e-9 W=180e-9 AD=18.9e-15 AS=18.9e-15 PD=390e-9 PS=390e-9 M=1
m0 out a net16 0 NMOS_VTL L=50e-9 W=180e-9 AD=18.9e-15 AS=18.9e-15 PD=390e-9 PS=390e-9 M=1
m3 out b vdd! vdd! PMOS_VTL L=50e-9 W=180e-9 AD=18.9e-15 AS=18.9e-15 PD=390e-9 PS=390e-9 M=1
m2 out a vdd! vdd! PMOS_VTL L=50e-9 W=180e-9 AD=18.9e-15 AS=18.9e-15 PD=390e-9 PS=390e-9 M=1
.ends NAND2
** End of subcircuit definition.

** Library name: my
** Cell name: AND2
** View name: schematic
.subckt AND2 a b out
xi0 net7 out INV
xi1 a b net7 NAND2
.ends AND2
** End of subcircuit definition.

** Library name: my
** Cell name: PC_CTRL
** View name: schematic
.subckt PC_CTRL _net1 _net0 a a_ b b_ pc
xi1 b net17 INV
xi0 a net18 INV
xi5 pc net17 _net0 AND2
xi4 pc b b_ AND2
xi3 a pc a_ AND2
xi2 net18 pc _net1 AND2
.ends PC_CTRL
** End of subcircuit definition.


.INCLUDE "MULT_TOP_v2.pex.netlist"

** Library name: my
** Cell name: MULT_TOP_v2_test
** View name: schematic
c31 s12 0 1e-15
c32 ov 0 1e-15
c3 s28 0 1e-15
c5 s26 0 1e-15
c4 s27 0 1e-15
c2 s29 0 1e-15
c8 s16 0 1e-15
c7 s24 0 1e-15
c10 s18 0 1e-15
c9 s17 0 1e-15
c6 s25 0 1e-15
c13 s22 0 1e-15
c12 s23 0 1e-15
c11 s19 0 1e-15
c16 s4 0 1e-15
c15 s20 0 1e-15
c18 s6 0 1e-15
c17 s5 0 1e-15
c14 s21 0 1e-15
c20 s3 0 1e-15
c21 s2 0 1e-15
c19 s7 0 1e-15
c23 s0 0 1e-15
c24 s8 0 1e-15
c25 s9 0 1e-15
c26 s10 0 1e-15
c22 s1 0 1e-15
c1 s30 0 1e-15
c0 s31 0 1e-15
c29 s14 0 1e-15
c27 s11 0 1e-15
c28 s15 0 1e-15
c30 s13 0 1e-15
v0 vdd! 0 DC=1.1
xi433 x2_b x3_b _x2 x2 _x3 x3 pc PC_CTRL
xi434 x4_b x5_b _x4 x4 _x5 x5 pc PC_CTRL
xi435 x6_b x7_b _x6 x6 _x7 x7 pc PC_CTRL
xi436 x0_b x1_b _x0 x0 _x1 x1 pc PC_CTRL
xi429 x8_b x9_b _x8 x8 _x9 x9 pc PC_CTRL
xi430 x10_b x11_b _x10 x10 _x11 x11 pc PC_CTRL
xi431 x12_b x13_b _x12 x12 _x13 x13 pc PC_CTRL
xi432 x14_b x15_b _x14 x14 _x15 x15 pc PC_CTRL
xi440 vdd_pc 0 0 gnd_pc 0 0 pc PC_CTRL
xi404 y6_b y7_b _y6 y6 _y7 y7 pc PC_CTRL
xi403 y4_b y5_b _y4 y4 _y5 y5 pc PC_CTRL
xi402 y2_b y3_b _y2 y2 _y3 y3 pc PC_CTRL
xi401 y0_b y1_b _y0 y0 _y1 y1 pc PC_CTRL
xi400 y14_b y15_b _y14 y14 _y15 y15 pc PC_CTRL
xi399 y12_b y13_b _y12 y12 _y13 y13 pc PC_CTRL
xi398 y10_b y11_b _y10 y10 _y11 y11 pc PC_CTRL
xi397 y8_b y9_b _y8 y8 _y9 y9 pc PC_CTRL


v250 pc 0 PULSE 0 1.1 0 10e-12 10e-12 120E-9 200e-9

v218	_x0		0	PULSE	!X0_	X0_		0	1.00E-11	1.00E-11	130e-09	200E-09
v246	_x1		0	PULSE	!X1_	X1_		0	1.00E-11	1.00E-11	130e-09	200E-09
v243	_x2		0	PULSE	!X2_	X2_		0	1.00E-11	1.00E-11	130e-09	200E-09
v247	_x3		0	PULSE	!X3_	X3_		0	1.00E-11	1.00E-11	130e-09	200E-09
v244	_x4		0	PULSE	!X4_	X4_		0	1.00E-11	1.00E-11	130e-09	200E-09
v248	_x5		0	PULSE	!X5_	X5_		0	1.00E-11	1.00E-11	130e-09	200E-09
v245	_x6		0	PULSE	!X6_	X6_		0	1.00E-11	1.00E-11	130e-09	200E-09
v249	_x7		0	PULSE	!X7_	X7_		0	1.00E-11	1.00E-11	130e-09	200E-09
v235	_x8		0	PULSE	!X8_	X8_		0	1.00E-11	1.00E-11	130e-09	200E-09
v239	_x9		0	PULSE	!X9_	X9_		0	1.00E-11	1.00E-11	130e-09	200E-09
v236	_x10	0	PULSE	!X10_	X10_	0	1.00E-11	1.00E-11	130e-09	200E-09
v240	_x11	0	PULSE	!X11_	X11_	0	1.00E-11	1.00E-11	130e-09	200E-09
v237	_x12	0	PULSE	!X12_	X12_	0	1.00E-11	1.00E-11	130e-09	200E-09
v241	_x13	0	PULSE	!X13_	X13_	0	1.00E-11	1.00E-11	130e-09	200E-09
v238	_x14	0	PULSE	!X14_	X14_	0	1.00E-11	1.00E-11	130e-09	200E-09
v242	_x15	0	PULSE	!X15_	X15_	0	1.00E-11	1.00E-11	130e-09	200E-09


v210	_y0		0	PULSE	!Y0_	Y0_		0	1.00E-11	1.00E-11	130e-09	200E-09
v214	_y1		0	PULSE	!Y1_	Y1_		0	1.00E-11	1.00E-11	130e-09	200E-09
v211	_y2		0	PULSE	!Y2_	Y2_		0	1.00E-11	1.00E-11	130e-09	200E-09
v215	_y3		0	PULSE	!Y3_	Y3_		0	1.00E-11	1.00E-11	130e-09	200E-09
v212	_y4		0	PULSE	!Y4_	Y4_		0	1.00E-11	1.00E-11	130e-09	200E-09
v216	_y5		0	PULSE	!Y5_	Y5_		0	1.00E-11	1.00E-11	130e-09	200E-09
v213	_y6		0	PULSE	!Y6_	Y6_		0	1.00E-11	1.00E-11	130e-09	200E-09
v217	_y7		0	PULSE	!Y7_	Y7_		0	1.00E-11	1.00E-11	130e-09	200E-09
v202	_y8		0	PULSE	!Y8_	Y8_		0	1.00E-11	1.00E-11	130e-09	200E-09
v206	_y9		0	PULSE	!Y9_	Y9_		0	1.00E-11	1.00E-11	130e-09	200E-09
v203	_y10	0	PULSE	!Y10_	Y10_	0	1.00E-11	1.00E-11	130e-09	200E-09
v207	_y11	0	PULSE	!Y11_	Y11_	0	1.00E-11	1.00E-11	130e-09	200E-09
v204	_y12	0	PULSE	!Y12_	Y12_	0	1.00E-11	1.00E-11	130e-09	200E-09
v208	_y13	0	PULSE	!Y13_	Y13_	0	1.00E-11	1.00E-11	130e-09	200E-09
v205	_y14	0	PULSE	!Y14_	Y14_	0	1.00E-11	1.00E-11	130e-09	200E-09
v209	_y15	0	PULSE	!Y15_	Y15_	0	1.00E-11	1.00E-11	130e-09	200E-09

xi489 VDD! GND! X15_B X15 X14_B X14 X13_B X13 X12_B X12 X11_B X11
+ X10_B X10 X9_B X9 Y15 Y15_B X8_B X8 X7_B X7 X6_B X6 X5_B X5 X4_B X4 X3_B X3
+ X2_B X2 X1_B X1 X0_B X0 Y13_B Y13 Y11_B Y11 Y9_B Y9 Y7_B Y7 Y5_B Y5 Y3_B Y3
+ Y1_B Y1 VDD_PC GND_PC Y14_B Y14 Y12_B Y12 Y10_B Y10 Y8_B Y8 Y6_B Y6 Y4_B Y4
+ Y2_B Y2 Y0_B Y0 OV S31 S30 S29 S28 S27 S26 S25 S24 S23 S22 S21 S20 S19 S18 S17
+ S16 S15 S14 S13 S12 S11 S10 S9 S8 S7 S6 S5 S4 S3 S2 S1 S0 MULT_TOP_v2



.END
