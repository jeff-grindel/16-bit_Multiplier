** Generated for: hspiceD
** Generated on: Jun 11 20:43:30 2013
** Design library name: my
** Design cell name: PPA_test
** Design view name: schematic
.GLOBAL vdd!

.TRAN 1e-12 5E-9 START=0.0 SWEEP DATA=D
.DATA D
+	A0_	A1_	A2_	A3_	A4_	A5_	A6_	A7_	A8_	A9_	A10_	A11_	A12_	A13_	A14_	A15_	A16_	A17_	A18_	A19_	A20_	A21_	A22_	A23_	A24_	A25_	A26_	A27_	A28_	A29_	A30_	A31_	B0_	B1_	B2_	B3_	B4_	B5_	B6_	B7_	B8_	B9_	B10_	B11_	B12_	B13_	B14_	B15_	B16_	B17_	B18_	B19_	B20_	B21_	B22_	B23_	B24_	B25_	B26_	B27_	B28_	B29_	B30_	B31_	!A0_	!A1_	!A2_	!A3_	!A4_	!A5_	!A6_	!A7_	!A8_	!A9_	!A10_	!A11_	!A12_	!A13_	!A14_	!A15_	!A16_	!A17_	!A18_	!A19_	!A20_	!A21_	!A22_	!A23_	!A24_	!A25_	!A26_	!A27_	!A28_	!A29_	!A30_	!A31_	!B0_	!B1_	!B2_	!B3_	!B4_	!B5_	!B6_	!B7_	!B8_	!B9_	!B10_	!B11_	!B12_	!B13_	!B14_	!B15_	!B16_	!B17_	!B18_	!B19_	!B20_	!B21_	!B22_	!B23_	!B24_	!B25_	!B26_	!B27_	!B28_	!B29_	!B30_	!B31_
**+	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1
**+	1.1	0	0	1.1	0	0	1.1	0	0	1.1	1.1	0	0	1.1	1.1	1.1	0	0	1.1	1.1	1.1	1.1	1.1	0	1.1	0	1.1	1.1	1.1	1.1	1.1	0	0	0	1.1	0	0	1.1	0	0	0	0	1.1	0	1.1	1.1	0	0	0	0	1.1	0	1.1	0	0	0	1.1	0	1.1	0	0	0	0	0	0	1.1	1.1	0	1.1	1.1	0	1.1	1.1	0	0	1.1	1.1	0	0	0	1.1	1.1	0	0	0	0	0	1.1	0	1.1	0	0	0	0	0	1.1	1.1	1.1	0	1.1	1.1	0	1.1	1.1	1.1	1.1	0	1.1	0	0	1.1	1.1	1.1	1.1	0	1.1	0	1.1	1.1	1.1	0	1.1	0	1.1	1.1	1.1	1.1	1.1
**+	1.1	0	1.1	1.1	1.1	0	1.1	0	0	0	0	1.1	0	0	0	1.1	1.1	0	0	1.1	1.1	1.1	1.1	1.1	1.1	1.1	0	1.1	1.1	0	1.1	1.1	1.1	1.1	0	1.1	1.1	1.1	1.1	0	1.1	0	0	1.1	1.1	0	0	0	1.1	0	1.1	1.1	0	1.1	0	0	0	1.1	0	1.1	0	0	0	0	0	1.1	0	0	0	1.1	0	1.1	1.1	1.1	1.1	0	1.1	1.1	1.1	0	0	1.1	1.1	0	0	0	0	0	0	0	1.1	0	0	1.1	0	0	0	0	1.1	0	0	0	0	1.1	0	1.1	1.1	0	0	1.1	1.1	1.1	0	1.1	0	0	1.1	0	1.1	1.1	1.1	0	1.1	0	1.1	1.1	1.1	1.1
**+	0	1.1	0	0	1.1	1.1	1.1	0	0	1.1	0	0	0	1.1	1.1	0	1.1	0	0	0	1.1	1.1	1.1	1.1	1.1	1.1	1.1	0	1.1	1.1	1.1	0	1.1	0	1.1	1.1	1.1	0	1.1	0	0	0	1.1	1.1	1.1	1.1	0	1.1	0	0	0	1.1	1.1	1.1	0	0	1.1	1.1	1.1	0	0	0	0	0	1.1	0	1.1	1.1	0	0	0	1.1	1.1	0	1.1	1.1	1.1	0	0	1.1	0	1.1	1.1	1.1	0	0	0	0	0	0	0	1.1	0	0	0	1.1	0	1.1	0	0	0	1.1	0	1.1	1.1	1.1	0	0	0	0	1.1	0	1.1	1.1	1.1	0	0	0	1.1	1.1	0	0	0	1.1	1.1	1.1	1.1	1.1
**+	0	1.1	1.1	1.1	1.1	0	1.1	1.1	1.1	1.1	0	0	0	1.1	0	0	0	1.1	1.1	1.1	0	1.1	1.1	1.1	1.1	0	0	1.1	0	1.1	0	0	1.1	0	1.1	1.1	1.1	1.1	0	0	1.1	0	0	0	1.1	1.1	0	0	1.1	0	1.1	0	0	0	0	1.1	0	0	1.1	1.1	0	0	1.1	1.1	1.1	0	0	0	0	1.1	0	0	0	0	1.1	1.1	1.1	0	1.1	1.1	1.1	0	0	0	1.1	0	0	0	0	1.1	1.1	0	1.1	0	1.1	1.1	0	1.1	0	0	0	0	1.1	1.1	0	1.1	1.1	1.1	0	0	1.1	1.1	0	1.1	0	1.1	1.1	1.1	1.1	0	1.1	1.1	0	0	1.1	1.1	0	0
**+	0	1.1	1.1	0	0	1.1	0	0	1.1	0	0	1.1	0	1.1	1.1	0	0	1.1	1.1	0	1.1	0	1.1	0	1.1	1.1	1.1	0	0	1.1	1.1	0	1.1	0	0	0	0	0	1.1	1.1	0	1.1	0	0	1.1	0	0	0	0	1.1	0	0	0	0	0	0	1.1	1.1	0	1.1	0	1.1	0	1.1	1.1	0	0	1.1	1.1	0	1.1	1.1	0	1.1	1.1	0	1.1	0	0	1.1	1.1	0	0	1.1	0	1.1	0	1.1	0	0	0	1.1	1.1	0	0	1.1	0	1.1	1.1	1.1	1.1	1.1	0	0	1.1	0	1.1	1.1	0	1.1	1.1	1.1	1.1	0	1.1	1.1	1.1	1.1	1.1	1.1	0	0	1.1	0	1.1	0	1.1	0
**+	1.1	1.1	0	1.1	0	1.1	1.1	0	1.1	0	0	1.1	1.1	0	0	1.1	1.1	0	1.1	0	1.1	0	1.1	0	0	0	1.1	1.1	1.1	0	0	1.1	1.1	0	1.1	0	1.1	1.1	0	0	0	0	0	1.1	0	0	0	0	1.1	1.1	1.1	0	0	1.1	0	1.1	0	0	1.1	1.1	1.1	1.1	1.1	1.1	0	0	1.1	0	1.1	0	0	1.1	0	1.1	1.1	0	0	1.1	1.1	0	0	1.1	0	1.1	0	1.1	0	1.1	1.1	1.1	0	0	0	1.1	1.1	0	0	1.1	0	1.1	0	0	1.1	1.1	1.1	1.1	1.1	0	1.1	1.1	1.1	1.1	0	0	0	1.1	1.1	0	1.1	0	1.1	1.1	0	0	0	0	0	0
**+	1.1	1.1	0	1.1	1.1	1.1	0	1.1	0	1.1	1.1	1.1	0	0	1.1	1.1	1.1	0	1.1	0	0	0	0	1.1	0	0	0	0	1.1	1.1	0	0	1.1	0	0	0	0	0	0	1.1	1.1	1.1	0	0	0	0	0	1.1	1.1	1.1	0	1.1	1.1	1.1	0	1.1	0	0	1.1	1.1	0	0	0	1.1	0	0	1.1	0	0	0	1.1	0	1.1	0	0	0	1.1	1.1	0	0	0	1.1	0	1.1	1.1	1.1	1.1	0	1.1	1.1	1.1	1.1	0	0	1.1	1.1	0	1.1	1.1	1.1	1.1	1.1	1.1	0	0	0	1.1	1.1	1.1	1.1	1.1	0	0	0	1.1	0	0	0	1.1	0	1.1	1.1	0	0	1.1	1.1	1.1	0
**+	0	0	0	1.1	1.1	0	1.1	0	1.1	1.1	0	1.1	0	1.1	0	1.1	0	1.1	1.1	1.1	0	0	1.1	1.1	0	0	1.1	1.1	1.1	0	1.1	0	0	1.1	0	1.1	1.1	1.1	0	1.1	0	0	0	0	0	0	1.1	0	1.1	0	0	1.1	1.1	1.1	0	1.1	1.1	0	0	1.1	0	1.1	0	1.1	1.1	1.1	1.1	0	0	1.1	0	1.1	0	0	1.1	0	1.1	0	1.1	0	1.1	0	0	0	1.1	1.1	0	0	1.1	1.1	0	0	0	1.1	0	1.1	1.1	0	1.1	0	0	0	1.1	0	1.1	1.1	1.1	1.1	1.1	1.1	0	1.1	0	1.1	1.1	0	0	0	1.1	0	0	1.1	1.1	0	1.1	0	1.1	0
+	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0
+	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1	1.1

.ENDDATA 

.OP

.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
+    POST
.INCLUDE "/apps/FreePDK45/ncsu_basekit/models/hspice/hspice_nom.include"

.PRINT TRAN POWER
.MEASURE TRAN avgpwr AVG POWER FROM 0 to 5e-9

** Library name: my
** Cell name: INV
** View name: schematic
.subckt INV in out
m0 out in vdd! vdd! PMOS_VTL L=50e-9 W=180e-9 AD=18.9e-15 AS=18.9e-15 PD=390e-9 PS=390e-9 M=1
m1 out in 0 0 NMOS_VTL L=50e-9 W=90e-9 AD=9.45e-15 AS=9.45e-15 PD=300e-9 PS=300e-9 M=1
.ends INV
** End of subcircuit definition.

** Library name: my
** Cell name: NAND2
** View name: schematic
.subckt NAND2 a b out
m1 net16 b 0 0 NMOS_VTL L=50e-9 W=180e-9 AD=18.9e-15 AS=18.9e-15 PD=390e-9 PS=390e-9 M=1
m0 out a net16 0 NMOS_VTL L=50e-9 W=180e-9 AD=18.9e-15 AS=18.9e-15 PD=390e-9 PS=390e-9 M=1
m3 out b vdd! vdd! PMOS_VTL L=50e-9 W=180e-9 AD=18.9e-15 AS=18.9e-15 PD=390e-9 PS=390e-9 M=1
m2 out a vdd! vdd! PMOS_VTL L=50e-9 W=180e-9 AD=18.9e-15 AS=18.9e-15 PD=390e-9 PS=390e-9 M=1
.ends NAND2
** End of subcircuit definition.

** Library name: my
** Cell name: AND2
** View name: schematic
.subckt AND2 a b out
xi0 net7 out INV
xi1 a b net7 NAND2
.ends AND2
** End of subcircuit definition.

** Library name: my
** Cell name: PC_CTRL
** View name: schematic
.subckt PC_CTRL _net1 _net0 a a_ b b_ pc
xi1 b net17 INV
xi0 a net18 INV
xi5 pc net17 _net0 AND2
xi4 pc b b_ AND2
xi3 a pc a_ AND2
xi2 net18 pc _net1 AND2
.ends PC_CTRL
** End of subcircuit definition.

.INCLUDE "PPA.pex.netlist"

** Library name: my
** Cell name: PPA_test
** View name: schematic
c32 ov 0 5e-15
c31 s24 0 1e-15
c30 s25 0 1e-15
c29 s26 0 1e-15
c28 s27 0 1e-15
c27 s20 0 1e-15
c26 s21 0 1e-15
c25 s22 0 1e-15
c24 s23 0 1e-15
c23 s16 0 1e-15
c22 s17 0 1e-15
c21 s18 0 1e-15
c20 s19 0 1e-15
c19 s12 0 1e-15
c18 s13 0 1e-15
c17 s14 0 1e-15
c16 s15 0 1e-15
c15 s11 0 1e-15
c14 s10 0 1e-15
c13 s9 0 1e-15
c12 s8 0 1e-15
c11 s7 0 1e-15
c10 s6 0 1e-15
c9 s5 0 1e-15
c8 s4 0 1e-15
c7 s28 0 1e-15
c6 s29 0 1e-15
c5 s30 0 1e-15
c4 s31 0 1e-15
c3 s0 0 1e-15
c2 s1 0 1e-15
c1 s2 0 1e-15
c0 s3 0 1e-15
v0 vdd! 0 DC=1.1
xi135 b16_b b17_b _b16 b16 _b17 b17 pc PC_CTRL
xi134 b18_b b19_b _b18 b18 _b19 b19 pc PC_CTRL
xi133 b20_b b21_b _b20 b20 _b21 b21 pc PC_CTRL
xi132 b22_b b23_b _b22 b22 _b23 b23 pc PC_CTRL
xi131 b26_b b27_b _b26 b26 _b27 b27 pc PC_CTRL
xi130 b28_b b29_b _b28 b28 _b29 b29 pc PC_CTRL
xi129 b30_b b31_b _b30 b30 _b31 b31 pc PC_CTRL
xi128 b24_b b25_b _b24 b24 _b25 b25 pc PC_CTRL
xi116 b6_b b7_b _b6 b6 _b7 b7 pc PC_CTRL
xi119 b4_b b5_b _b4 b4 _b5 b5 pc PC_CTRL
xi118 b2_b b3_b _b2 b2 _b3 b3 pc PC_CTRL
xi117 b0_b b1_b _b0 b0 _b1 b1 pc PC_CTRL
xi103 a26_b a27_b _a26 a26 _a27 a27 pc PC_CTRL
xi102 a28_b a29_b _a28 a28 _a29 a29 pc PC_CTRL
xi101 a30_b a31_b _a30 a30 _a31 a31 pc PC_CTRL
xi100 a24_b a25_b _a24 a24 _a25 a25 pc PC_CTRL
xi95 a18_b a19_b _a18 a18 _a19 a19 pc PC_CTRL
xi94 a20_b a21_b _a20 a20 _a21 a21 pc PC_CTRL
xi93 a22_b a23_b _a22 a22 _a23 a23 pc PC_CTRL
xi92 a16_b a17_b _a16 a16 _a17 a17 pc PC_CTRL
xi87 a10_b a11_b _a10 a10 _a11 a11 pc PC_CTRL
xi86 a12_b a13_b _a12 a12 _a13 a13 pc PC_CTRL
xi85 a14_b a15_b _a14 a14 _a15 a15 pc PC_CTRL
xi84 a8_b a9_b _a8 a8 _a9 a9 pc PC_CTRL
xi70 b8_b b9_b _b8 b8 _b9 b9 pc PC_CTRL
xi68 b10_b b11_b _b10 b10 _b11 b11 pc PC_CTRL
xi66 b12_b b13_b _b12 b12 _b13 b13 pc PC_CTRL
xi64 b14_b b15_b _b14 b14 _b15 b15 pc PC_CTRL
xi79 a2_b a3_b _a2 a2 _a3 a3 pc PC_CTRL
xi77 a6_b a7_b _a6 a6 _a7 a7 pc PC_CTRL
xi78 a4_b a5_b _a4 a4 _a5 a5 pc PC_CTRL
xi76 a0_b a1_b _a0 a0 _a1 a1 pc PC_CTRL

v26	_a0	0	PULSE	!A0_	A0_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v31	_a1	0	PULSE	!A1_	A1_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v25	_a2	0	PULSE	!A2_	A2_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v30	_a3	0	PULSE	!A3_	A3_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v24	_a4	0	PULSE	!A4_	A4_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v29	_a5	0	PULSE	!A5_	A5_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v27	_a6	0	PULSE	!A6_	A6_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v28	_a7	0	PULSE	!A7_	A7_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v34	_a8	0	PULSE	!A8_	A8_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v39	_a9	0	PULSE	!A9_	A9_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v33	_a10	0	PULSE	!A10_	A10_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v38	_a11	0	PULSE	!A11_	A11_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v32	_a12	0	PULSE	!A12_	A12_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v37	_a13	0	PULSE	!A13_	A13_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v35	_a14	0	PULSE	!A14_	A14_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v36	_a15	0	PULSE	!A15_	A15_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v42	_a16	0	PULSE	!A16_	A16_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v47	_a17	0	PULSE	!A17_	A17_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v41	_a18	0	PULSE	!A18_	A18_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v46	_a19	0	PULSE	!A19_	A19_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v40	_a20	0	PULSE	!A20_	A20_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v45	_a21	0	PULSE	!A21_	A21_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v43	_a22	0	PULSE	!A22_	A22_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v44	_a23	0	PULSE	!A23_	A23_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v50	_a24	0	PULSE	!A24_	A24_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v55	_a25	0	PULSE	!A25_	A25_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v49	_a26	0	PULSE	!A26_	A26_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v54	_a27	0	PULSE	!A27_	A27_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v48	_a28	0	PULSE	!A28_	A28_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v53	_a29	0	PULSE	!A29_	A29_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v51	_a30	0	PULSE	!A30_	A30_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v52	_a31	0	PULSE	!A31_	A31_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09





v65	_b0	0	PULSE	!B0_	B0_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v69	_b1	0	PULSE	!B1_	B1_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v64	_b2	0	PULSE	!B2_	B2_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v68	_b3	0	PULSE	!B3_	B3_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v66	_b4	0	PULSE	!B4_	B4_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v70	_b5	0	PULSE	!B5_	B5_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v67	_b6	0	PULSE	!B6_	B6_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v71	_b7	0	PULSE	!B7_	B7_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v23	_b8	0	PULSE	!B8_	B8_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v22	_b9	0	PULSE	!B9_	B9_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v21	_b10	0	PULSE	!B10_	B10_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v20	_b11	0	PULSE	!B11_	B11_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v19	_b12	0	PULSE	!B12_	B12_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v18	_b13	0	PULSE	!B13_	B13_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v17	_b14	0	PULSE	!B14_	B14_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v16	_b15	0	PULSE	!B15_	B15_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v81	_b16	0	PULSE	!B16_	B16_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v86	_b17	0	PULSE	!B17_	B17_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v82	_b18	0	PULSE	!B18_	B18_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v87	_b19	0	PULSE	!B19_	B19_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v80	_b20	0	PULSE	!B20_	B20_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v85	_b21	0	PULSE	!B21_	B21_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v83	_b22	0	PULSE	!B22_	B22_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v84	_b23	0	PULSE	!B23_	B23_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v74	_b24	0	PULSE	!B24_	B24_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v79	_b25	0	PULSE	!B25_	B25_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v73	_b26	0	PULSE	!B26_	B26_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v78	_b27	0	PULSE	!B27_	B27_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v72	_b28	0	PULSE	!B28_	B28_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v77	_b29	0	PULSE	!B29_	B29_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v75	_b30	0	PULSE	!B30_	B30_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09
v76	_b31	0	PULSE	!B31_	B31_	0.00E+00	1.00E-11	1.00E-11	3.00E-09	5.00E-09


v1 pc 0 PULSE 0 1.1 0 10e-12 10e-12 2.6E-9 5E-9

xi34 OV GND! VDD! S31 A31 A31_B B31 B31_B S30 A30 A30_B B30 B30_B S29
+ A29 A29_B B29 B29_B S28 A28 A28_B B28 B28_B S27 A27 A27_B B27 B27_B S26 A26
+ A26_B B26 B26_B S25 A25 A25_B B25 B25_B S24 A24 A24_B B24 B24_B S23 A23 A23_B
+ B23 B23_B S22 A22 A22_B B22 B22_B S21 A21 A21_B B21 B21_B S20 A20 A20_B B20
+ B20_B S19 A19 A19_B B19 B19_B S18 A18 A18_B B18 B18_B S17 A17 A17_B B17 B17_B
+ S16 A16 A16_B B16 B16_B S15 A15 A15_B B15 B15_B S14 A14 A14_B B14 B14_B S13
+ A13 A13_B B13 B13_B S12 A12 A12_B B12 B12_B S11 A11 A11_B B11 B11_B S10 A10
+ A10_B B10 B10_B S9 A9 A9_B B9 B9_B S8 A8 A8_B B8 B8_B S7 A7 A7_B B7 B7_B S6 A6
+ A6_B B6 B6_B S5 A5 A5_B B5 B5_B S4 A4 A4_B B4 B4_B S3 A3 A3_B B3 B3_B S2 A2
+ A2_B B2 B2_B S1 A1 A1_B B1 B1_B S0 A0 A0_B B0 B0_B PPA
.END
