* SPICE NETLIST
***************************************

.SUBCKT NAND2 a gnd! b OUT vdd!
** N=6 EP=5 IP=0 FDC=4
M0 6 a gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07 $X=210 $Y=-360 $D=1
M1 OUT b 6 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=2.52e-14 PD=5.75e-07 PS=6.4e-07 $X=590 $Y=-360 $D=1
M2 OUT a vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07 $X=210 $Y=670 $D=0
M3 vdd! b OUT vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14 PD=5.7e-07 PS=6.4e-07 $X=590 $Y=670 $D=0
.ENDS
***************************************
.SUBCKT SP_XOR_DR A P !A !P B gnd! vdd! !B
** N=14 EP=8 IP=10 FDC=22
M0 1 !B gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.025e-14 PD=6.4e-07 PS=5.85e-07 $X=675 $Y=110 $D=1
M1 3 A 1 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=2.52e-14 PD=6.65e-07 PS=6.4e-07 $X=1055 $Y=110 $D=1
M2 6 !A 1 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=5.445e-14 PD=6.65e-07 PS=9.65e-07 $X=2685 $Y=110 $D=1
M3 9 B gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.025e-14 PD=6.4e-07 PS=5.85e-07 $X=3955 $Y=110 $D=1
M4 10 !A 9 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=2.52e-14 PD=6.65e-07 PS=6.4e-07 $X=4335 $Y=110 $D=1
M5 14 A 9 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=5.445e-14 PD=6.65e-07 PS=9.65e-07 $X=5965 $Y=110 $D=1
M6 3 A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=675 $Y=3505 $D=0
M7 vdd! P 3 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=1495 $Y=3505 $D=0
M8 6 !A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=2305 $Y=3505 $D=0
M9 vdd! !P 6 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3125 $Y=3505 $D=0
M10 10 !A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=3955 $Y=3505 $D=0
M11 vdd! P 10 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=4775 $Y=3505 $D=0
M12 14 A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=5585 $Y=3505 $D=0
M13 vdd! !P 14 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=6405 $Y=3505 $D=0
X14 14 gnd! 6 !P vdd! NAND2 $T=7820 250 0 0 $X=7370 $Y=-395
X15 3 gnd! 10 P vdd! NAND2 $T=7820 3040 0 0 $X=7370 $Y=2395
.ENDS
***************************************
