* SPICE NETLIST
***************************************

.SUBCKT NAND2 A gnd! B OUT vdd!
** N=6 EP=5 IP=0 FDC=4
M0 6 A gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07 $X=210 $Y=-360 $D=1
M1 OUT B 6 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=2.52e-14 PD=5.75e-07 PS=6.4e-07 $X=590 $Y=-360 $D=1
M2 OUT A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07 $X=210 $Y=670 $D=0
M3 vdd! B OUT vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14 PD=5.7e-07 PS=6.4e-07 $X=590 $Y=670 $D=0
.ENDS
***************************************
.SUBCKT SP_XOR3_DR C_b B_b A A_b B P C P_b gnd! vdd!
** N=20 EP=10 IP=10 FDC=28
M0 17 C_b gnd! gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=4.995e-14 AS=3.0375e-14 PD=9.1e-07 PS=7.65e-07 $X=-545 $Y=-1090 $D=1
M1 4 B_b 17 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=5.1975e-14 AS=4.995e-14 PD=9.25e-07 PS=9.1e-07 $X=-75 $Y=-1090 $D=1
M2 18 B 4 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=4.7925e-14 AS=5.1975e-14 PD=8.95e-07 PS=9.25e-07 $X=410 $Y=-1090 $D=1
M3 gnd! C 18 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=3.4425e-14 AS=4.7925e-14 PD=7.95e-07 PS=8.95e-07 $X=865 $Y=-1090 $D=1
M4 4 A 7 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=5.6025e-14 AS=4.185e-14 PD=9.55e-07 PS=8.5e-07 $X=1790 $Y=-1090 $D=1
M5 10 A_b 4 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=4.1175e-14 AS=5.6025e-14 PD=8.45e-07 PS=9.55e-07 $X=2305 $Y=-1090 $D=1
M6 19 C gnd! gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=4.995e-14 AS=3.0375e-14 PD=9.1e-07 PS=7.65e-07 $X=3485 $Y=-1090 $D=1
M7 12 B_b 19 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=5.1975e-14 AS=4.995e-14 PD=9.25e-07 PS=9.1e-07 $X=3955 $Y=-1090 $D=1
M8 20 B 12 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=4.7925e-14 AS=5.1975e-14 PD=8.95e-07 PS=9.25e-07 $X=4440 $Y=-1090 $D=1
M9 gnd! C_b 20 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=3.4425e-14 AS=4.7925e-14 PD=7.95e-07 PS=8.95e-07 $X=4895 $Y=-1090 $D=1
M10 12 A_b 13 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=5.6025e-14 AS=4.185e-14 PD=9.55e-07 PS=8.5e-07 $X=5820 $Y=-1090 $D=1
M11 16 A 12 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=4.1175e-14 AS=5.6025e-14 PD=8.45e-07 PS=9.55e-07 $X=6335 $Y=-1090 $D=1
M12 7 A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=-30 $Y=4245 $D=0
M13 vdd! P 7 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=790 $Y=4245 $D=0
M14 10 A_b vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=2305 $Y=4245 $D=0
M15 vdd! P_b 10 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3125 $Y=4245 $D=0
M16 13 A_b vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=3955 $Y=4245 $D=0
M17 vdd! P 13 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=4775 $Y=4245 $D=0
M18 16 A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=6335 $Y=4245 $D=0
M19 vdd! P_b 16 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=7155 $Y=4245 $D=0
X20 16 gnd! 10 P_b vdd! NAND2 $T=9525 -770 0 0 $X=9075 $Y=-1415
X21 7 gnd! 13 P vdd! NAND2 $T=9525 3780 0 0 $X=9075 $Y=3135
.ENDS
***************************************
