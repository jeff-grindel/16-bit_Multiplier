* SPICE NETLIST
***************************************

.SUBCKT M2_M1_via
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT NAND2 A gnd! B OUT vdd!
** N=6 EP=5 IP=0 FDC=4
M0 6 A gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07 $X=210 $Y=-360 $D=1
M1 OUT B 6 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=2.52e-14 PD=5.75e-07 PS=6.4e-07 $X=590 $Y=-360 $D=1
M2 OUT A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07 $X=210 $Y=670 $D=0
M3 vdd! B OUT vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14 PD=5.7e-07 PS=6.4e-07 $X=590 $Y=670 $D=0
.ENDS
***************************************
.SUBCKT SP_MAJ IN0 IN1 IN2 OUT gnd! vdd!
** N=10 EP=6 IP=5 FDC=13
M0 7 IN1 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.025e-14 PD=6.4e-07 PS=5.85e-07 $X=675 $Y=-190 $D=1
M1 gnd! IN2 7 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=2.52e-14 PD=6.65e-07 PS=6.4e-07 $X=1055 $Y=-190 $D=1
M2 5 IN0 7 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.115e-14 PD=5.85e-07 PS=5.95e-07 $X=1925 $Y=-190 $D=1
M3 10 IN2 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.745e-14 PD=6.4e-07 PS=6.65e-07 $X=2745 $Y=-190 $D=1
M4 6 IN1 10 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.52e-14 PD=5.85e-07 PS=6.4e-07 $X=3125 $Y=-190 $D=1
M5 5 IN0 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=675 $Y=2740 $D=0
M6 vdd! OUT 5 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=1495 $Y=2740 $D=0
M7 6 OUT vdd! vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=2305 $Y=2740 $D=0
M8 vdd! IN1 6 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=3125 $Y=2740 $D=0
X9 5 gnd! 6 OUT vdd! NAND2 $T=4925 170 0 0 $X=4475 $Y=-475
.ENDS
***************************************
.SUBCKT SP_FA_DR vdd! A B C A_b gnd! B_b C_b S S_b Co Co_b
** N=22 EP=12 IP=28 FDC=54
M0 14 A 18 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=5.6025e-14 AS=4.1175e-14 PD=9.55e-07 PS=8.45e-07 $X=19835 $Y=6770 $D=1
M1 9 A_b 14 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=4.185e-14 AS=5.6025e-14 PD=8.5e-07 PS=9.55e-07 $X=19835 $Y=7285 $D=1
M2 19 C_b gnd! gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=4.7925e-14 AS=3.4425e-14 PD=8.95e-07 PS=7.95e-07 $X=19835 $Y=8210 $D=1
M3 14 B 19 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=5.1975e-14 AS=4.7925e-14 PD=9.25e-07 PS=8.95e-07 $X=19835 $Y=8665 $D=1
M4 20 B_b 14 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=4.995e-14 AS=5.1975e-14 PD=9.1e-07 PS=9.25e-07 $X=19835 $Y=9150 $D=1
M5 gnd! C 20 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=3.0375e-14 AS=4.995e-14 PD=7.65e-07 PS=9.1e-07 $X=19835 $Y=9620 $D=1
M6 15 A_b 13 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=5.6025e-14 AS=4.1175e-14 PD=9.55e-07 PS=8.45e-07 $X=19835 $Y=10800 $D=1
M7 11 A 15 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=4.185e-14 AS=5.6025e-14 PD=8.5e-07 PS=9.55e-07 $X=19835 $Y=11315 $D=1
M8 21 C gnd! gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=4.7925e-14 AS=3.4425e-14 PD=8.95e-07 PS=7.95e-07 $X=19835 $Y=12240 $D=1
M9 15 B 21 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=5.1975e-14 AS=4.7925e-14 PD=9.25e-07 PS=8.95e-07 $X=19835 $Y=12695 $D=1
M10 22 B_b 15 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=4.995e-14 AS=5.1975e-14 PD=9.1e-07 PS=9.25e-07 $X=19835 $Y=13180 $D=1
M11 gnd! C_b 22 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=3.0375e-14 AS=4.995e-14 PD=7.65e-07 PS=9.1e-07 $X=19835 $Y=13650 $D=1
M12 vdd! A 18 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=14680 $Y=6770 $D=0
M13 vdd! A_b 9 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=14680 $Y=9150 $D=0
M14 vdd! A_b 13 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=14680 $Y=10800 $D=0
M15 vdd! A 11 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=14680 $Y=13135 $D=0
M16 18 S_b vdd! vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=14860 $Y=5950 $D=0
M17 9 S vdd! vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=14860 $Y=8330 $D=0
M18 13 S_b vdd! vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=14860 $Y=9980 $D=0
M19 11 S vdd! vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=14860 $Y=12315 $D=0
X26 11 gnd! 9 S vdd! NAND2 $T=15505 3680 1 270 $X=14175 $Y=2665
X27 18 gnd! 13 S_b vdd! NAND2 $T=20055 3680 1 270 $X=18725 $Y=2665
X28 A B C Co gnd! vdd! SP_MAJ $T=7925 12160 1 270 $X=4320 $Y=5760
X29 A_b B_b C_b Co_b gnd! vdd! SP_MAJ $T=12595 12160 1 270 $X=8990 $Y=5760
.ENDS
***************************************
.SUBCKT ICV_2
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT INV in gnd! vdd! out
** N=4 EP=4 IP=0 FDC=2
M0 out in gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07 $X=210 $Y=-180 $D=1
M1 out in vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07 $X=210 $Y=800 $D=0
.ENDS
***************************************
.SUBCKT SP_AND_DR out !A out_b !B gnd! vdd! B A
** N=12 EP=8 IP=9 FDC=16
M0 12 B gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.025e-14 PD=6.4e-07 PS=5.85e-07 $X=675 $Y=110 $D=1
M1 1 A 12 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=2.52e-14 PD=6.65e-07 PS=6.4e-07 $X=1055 $Y=110 $D=1
M2 4 !A gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=2305 $Y=110 $D=1
M3 11 !B gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3935 $Y=110 $D=1
M4 1 A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=675 $Y=3505 $D=0
M5 vdd! out 1 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=1495 $Y=3505 $D=0
M6 4 !A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=2305 $Y=3505 $D=0
M7 vdd! out_b 4 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3125 $Y=3505 $D=0
M8 11 !B vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=3935 $Y=3505 $D=0
M9 vdd! out_b 11 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=4755 $Y=3505 $D=0
X10 11 gnd! 4 out_b vdd! NAND2 $T=6255 250 0 0 $X=5805 $Y=-395
X11 1 gnd! vdd! out INV $T=6065 2910 0 0 $X=5615 $Y=2395
.ENDS
***************************************
.SUBCKT SP_OR_DR out_b A out B gnd! vdd! !B !A
** N=12 EP=8 IP=9 FDC=16
M0 12 !B gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.025e-14 PD=6.4e-07 PS=5.85e-07 $X=675 $Y=110 $D=1
M1 1 !A 12 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=2.52e-14 PD=6.65e-07 PS=6.4e-07 $X=1055 $Y=110 $D=1
M2 4 A gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=2305 $Y=110 $D=1
M3 11 B gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3935 $Y=110 $D=1
M4 1 !A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=675 $Y=3505 $D=0
M5 vdd! out_b 1 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=1495 $Y=3505 $D=0
M6 4 A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=2305 $Y=3505 $D=0
M7 vdd! out 4 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3125 $Y=3505 $D=0
M8 11 B vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=3935 $Y=3505 $D=0
M9 vdd! out 11 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=4755 $Y=3505 $D=0
X10 11 gnd! 4 out vdd! NAND2 $T=6255 250 0 0 $X=5805 $Y=-395
X11 1 gnd! vdd! out_b INV $T=6065 2910 0 0 $X=5615 $Y=2395
.ENDS
***************************************
.SUBCKT SP_XOR_DR A P !A !P B gnd! vdd! !B
** N=14 EP=8 IP=10 FDC=22
M0 1 !B gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.025e-14 PD=6.4e-07 PS=5.85e-07 $X=675 $Y=110 $D=1
M1 3 A 1 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=2.52e-14 PD=6.65e-07 PS=6.4e-07 $X=1055 $Y=110 $D=1
M2 6 !A 1 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=5.445e-14 PD=6.65e-07 PS=9.65e-07 $X=2685 $Y=110 $D=1
M3 9 B gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.025e-14 PD=6.4e-07 PS=5.85e-07 $X=3955 $Y=110 $D=1
M4 10 !A 9 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=2.52e-14 PD=6.65e-07 PS=6.4e-07 $X=4335 $Y=110 $D=1
M5 14 A 9 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=5.445e-14 PD=6.65e-07 PS=9.65e-07 $X=5965 $Y=110 $D=1
M6 3 A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=675 $Y=3505 $D=0
M7 vdd! P 3 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=1495 $Y=3505 $D=0
M8 6 !A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=2305 $Y=3505 $D=0
M9 vdd! !P 6 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3125 $Y=3505 $D=0
M10 10 !A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=3955 $Y=3505 $D=0
M11 vdd! P 10 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=4775 $Y=3505 $D=0
M12 14 A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=5585 $Y=3505 $D=0
M13 vdd! !P 14 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=6405 $Y=3505 $D=0
X14 14 gnd! 6 !P vdd! NAND2 $T=7820 250 0 0 $X=7370 $Y=-395
X15 3 gnd! 10 P vdd! NAND2 $T=7820 3040 0 0 $X=7370 $Y=2395
.ENDS
***************************************
.SUBCKT PPG_Cell_v1 POS_b POS TWO_b TWO Xj-1 Xj-1_b ONE_b Xj_b Xj vdd! PPG PPG_b ONE gnd!
** N=20 EP=14 IP=32 FDC=70
X0 11 TWO_b 12 Xj-1_b gnd! vdd! Xj-1 TWO SP_AND_DR $T=6270 10385 0 0 $X=6265 $Y=9990
X1 13 ONE_b 19 Xj_b gnd! vdd! Xj ONE SP_AND_DR $T=6270 16575 0 0 $X=6265 $Y=16180
X2 14 11 15 13 gnd! vdd! 19 12 SP_OR_DR $T=15980 16575 0 0 $X=15975 $Y=16180
X3 POS PPG POS_b PPG_b 15 gnd! vdd! 14 SP_XOR_DR $T=25595 16575 0 0 $X=25595 $Y=16180
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18
** N=18 EP=18 IP=28 FDC=140
X0 10 11 8 9 5 4 6 2 3 12 13 14 7 1 PPG_Cell_v1 $T=0 0 0 0 $X=1100 $Y=9990
X1 10 11 8 9 16 15 6 4 5 12 17 18 7 1 PPG_Cell_v1 $T=0 11630 0 0 $X=1100 $Y=21620
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26
** N=26 EP=26 IP=36 FDC=280
X0 1 2 3 11 12 4 5 6 7 8 9 10 15 16 13 14 17 18 ICV_3 $T=0 0 0 0 $X=1100 $Y=9990
X1 1 13 14 19 20 4 5 6 7 8 9 10 23 24 21 22 25 26 ICV_3 $T=0 23230 0 0 $X=1100 $Y=33220
.ENDS
***************************************
.SUBCKT PPG_Blk_v1 gnd! VDD_PC GND_PC PPGi_SE ONE_b ONE TWO_b TWO Yj+1_b PPGi_SE_b Yj+1 vdd! X15_b X15 PPGi+16 PPGi+16_b X14_b X14 PPGi+15 PPGi+15_b
+ X13_b X13 PPGi+14 PPGi+14_b X12_b X12 PPGi+13 PPGi+13_b X11_b X11 PPGi+12 PPGi+12_b X10_b X10 PPGi+11 PPGi+11_b X9_b X9 PPGi+10 PPGi+10_b
+ X8_b X8 PPGi+9 PPGi+9_b PPGi+8 PPGi+8_b PPGi+7 PPGi+7_b PPGi+6 PPGi+6_b PPGi+5 PPGi+5_b PPGi+4 PPGi+4_b PPGi+3 PPGi+3_b PPGi+2 PPGi+2_b PPGi+1 PPGi+1_b
+ X7_b PPGi PPGi_b X7 X6_b X6 X5_b X5 X4_b X4 X3_b X3 X2_b X2 X1_b X1 X0_b X0
** N=78 EP=78 IP=138 FDC=1260
X6 Yj+1_b Yj+1 TWO_b TWO GND_PC VDD_PC ONE_b VDD_PC GND_PC vdd! PPGi_SE PPGi_SE_b ONE gnd! PPG_Cell_v1 $T=23990 70620 0 270 $X=33980 $Y=32190
X7 Yj+1_b Yj+1 TWO_b TWO GND_PC VDD_PC ONE_b X0_b X0 vdd! PPGi PPGi_b ONE gnd! PPG_Cell_v1 $T=221505 70620 0 270 $X=231495 $Y=32190
X8 gnd! VDD_PC GND_PC ONE_b ONE TWO_b TWO Yj+1_b Yj+1 vdd! X15_b X15 X14_b X14 PPGi+16 PPGi+16_b PPGi+15 PPGi+15_b X13_b X13
+ X12_b X12 PPGi+14 PPGi+14_b PPGi+13 PPGi+13_b
+ ICV_4 $T=35625 70620 0 270 $X=45615 $Y=32190
X9 gnd! X12_b X12 ONE_b ONE TWO_b TWO Yj+1_b Yj+1 vdd! X11_b X11 X10_b X10 PPGi+12 PPGi+12_b PPGi+11 PPGi+11_b X9_b X9
+ X8_b X8 PPGi+10 PPGi+10_b PPGi+9 PPGi+9_b
+ ICV_4 $T=82095 70620 0 270 $X=92085 $Y=32190
X10 gnd! X8_b X8 ONE_b ONE TWO_b TWO Yj+1_b Yj+1 vdd! X7_b X7 X6_b X6 PPGi+8 PPGi+8_b PPGi+7 PPGi+7_b X5_b X5
+ X4_b X4 PPGi+6 PPGi+6_b PPGi+5 PPGi+5_b
+ ICV_4 $T=128565 70620 0 270 $X=138555 $Y=32190
X11 gnd! X4_b X4 ONE_b ONE TWO_b TWO Yj+1_b Yj+1 vdd! X3_b X3 X2_b X2 PPGi+4 PPGi+4_b PPGi+3 PPGi+3_b X1_b X1
+ X0_b X0 PPGi+2 PPGi+2_b PPGi+1 PPGi+1_b
+ ICV_4 $T=175035 70620 0 270 $X=185025 $Y=32190
.ENDS
***************************************
.SUBCKT PG_Blk !A A B !B gnd! vdd! !G G P !P
** N=10 EP=10 IP=16 FDC=38
X0 G !A !G !B gnd! vdd! B A SP_AND_DR $T=1500 3355 0 0 $X=1495 $Y=2960
X1 A P !A !P B gnd! vdd! !B SP_XOR_DR $T=1500 8640 0 0 $X=1500 $Y=8245
.ENDS
***************************************
.SUBCKT SP_XOR P !A B !B A gnd! vdd!
** N=11 EP=7 IP=5 FDC=12
M0 10 !B gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.025e-14 PD=6.4e-07 PS=5.85e-07 $X=675 $Y=110 $D=1
M1 1 A 10 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=2.52e-14 PD=6.65e-07 PS=6.4e-07 $X=1055 $Y=110 $D=1
M2 11 !A 3 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.745e-14 PD=6.4e-07 PS=6.65e-07 $X=2745 $Y=110 $D=1
M3 gnd! B 11 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.52e-14 PD=5.85e-07 PS=6.4e-07 $X=3125 $Y=110 $D=1
M4 1 A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=675 $Y=2740 $D=0
M5 vdd! P 1 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=1495 $Y=2740 $D=0
M6 3 P vdd! vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=2305 $Y=2740 $D=0
M7 vdd! !A 3 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=3125 $Y=2740 $D=0
X8 1 gnd! 3 P vdd! NAND2 $T=4925 470 0 0 $X=4475 $Y=-175
.ENDS
***************************************
.SUBCKT GREY_CELL !Gi-1 Gi-1 !Gi Gi !Pi Pi !G G gnd! vdd!
** N=15 EP=10 IP=9 FDC=18
M0 14 !Gi 7 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07 $X=1045 $Y=110 $D=1
M1 14 !Gi-1 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07 $X=1915 $Y=110 $D=1
M2 gnd! !Pi 14 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14 PD=5.7e-07 PS=6.4e-07 $X=2295 $Y=110 $D=1
M3 gnd! Gi 9 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3125 $Y=110 $D=1
M4 15 Gi-1 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.88e-14 AS=2.025e-14 PD=6.8e-07 PS=5.85e-07 $X=3935 $Y=110 $D=1
M5 11 Pi 15 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.385e-14 AS=2.88e-14 PD=6.25e-07 PS=6.8e-07 $X=4355 $Y=110 $D=1
M6 7 !Gi vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=675 $Y=3505 $D=0
M7 vdd! !G 7 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=1495 $Y=3505 $D=0
M8 9 Gi vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=2305 $Y=3505 $D=0
M9 vdd! G 9 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3125 $Y=3505 $D=0
M10 11 Pi vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=3935 $Y=3505 $D=0
M11 vdd! G 11 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=4755 $Y=3505 $D=0
X12 9 gnd! 11 G vdd! NAND2 $T=6185 3040 0 0 $X=5735 $Y=2395
X13 7 gnd! vdd! !G INV $T=6605 120 0 0 $X=6155 $Y=-395
.ENDS
***************************************
.SUBCKT BLACK_CELL Pi-1 !Pi-1 Gi !Gi Pi !Pi !Gi-1 gnd! vdd! Gi-1 !G G !P P
** N=14 EP=14 IP=18 FDC=34
X0 P !Pi !P !Pi-1 gnd! vdd! Pi-1 Pi SP_AND_DR $T=15 10675 0 0 $X=10 $Y=10280
X1 !Gi-1 Gi-1 !Gi Gi !Pi Pi !G G gnd! vdd! GREY_CELL $T=15 5615 0 0 $X=0 $Y=5220
.ENDS
***************************************
.SUBCKT PPA_v1 OV gnd! vdd! GND_PC S31 A31 A31_b B31 B31_b S30 A30 A30_b B30 B30_b S29 A29 A29_b B29 B29_b S28
+ A28 A28_b B28 B28_b S27 A27 A27_b B27 B27_b S26 A26 A26_b B26 B26_b S25 A25 A25_b B25 B25_b S24
+ A24 A24_b B24 B24_b S23 A23 A23_b B23 B23_b S22 A22 A22_b B22 B22_b S21 A21 A21_b B21 B21_b S20
+ A20 A20_b B20 B20_b S19 A19 A19_b B19 B19_b S18 A18 A18_b B18 B18_b S17 A17 A17_b B17 B17_b S16
+ A16 A16_b B16 B16_b S15 A15 A15_b B15 B15_b S14 A14 A14_b B14 B14_b S13 A13 A13_b B13 B13_b S12
+ A12 A12_b B12 B12_b S11 A11 A11_b B11 B11_b S10 A10 A10_b B10 B10_b S9 A9 A9_b B9 B9_b S8
+ A8 A8_b B8 B8_b S7 A7 A7_b B7 B7_b S6 A6 A6_b B6 B6_b S5 A5 A5_b B5 B5_b S4
+ A4 A4_b B4 B4_b S3 A3 A3_b B3 B3_b S2 A2 A2_b B2 B2_b S1 A1 A1_b B1 B1_b VDD_PC
+ S0 A0 A0_b B0 B0_b
** N=745 EP=165 IP=2226 FDC=5490
X0 A31_b A31 B31 B31_b gnd! vdd! 640 632 166 167 PG_Blk $T=-115700 210235 1 270 $X=-128710 $Y=198830
X1 A30_b A30 B30 B30_b gnd! vdd! 186 181 173 177 PG_Blk $T=-101650 210235 1 270 $X=-114660 $Y=198830
X2 A29_b A29 B29 B29_b gnd! vdd! 206 201 193 197 PG_Blk $T=-87600 210235 1 270 $X=-100610 $Y=198830
X3 A28_b A28 B28 B28_b gnd! vdd! 226 221 213 217 PG_Blk $T=-73550 210235 1 270 $X=-86560 $Y=198830
X4 A27_b A27 B27 B27_b gnd! vdd! 246 241 233 237 PG_Blk $T=-59500 210235 1 270 $X=-72510 $Y=198830
X5 A26_b A26 B26 B26_b gnd! vdd! 265 260 252 256 PG_Blk $T=-45450 210235 1 270 $X=-58460 $Y=198830
X6 A25_b A25 B25 B25_b gnd! vdd! 286 281 273 277 PG_Blk $T=-31400 210235 1 270 $X=-44410 $Y=198830
X7 A24_b A24 B24 B24_b gnd! vdd! 306 301 293 297 PG_Blk $T=-17350 210235 1 270 $X=-30360 $Y=198830
X8 A23_b A23 B23 B23_b gnd! vdd! 326 321 313 317 PG_Blk $T=-3300 210235 1 270 $X=-16310 $Y=198830
X9 A22_b A22 B22 B22_b gnd! vdd! 345 340 332 336 PG_Blk $T=10750 210235 1 270 $X=-2260 $Y=198830
X10 A21_b A21 B21 B21_b gnd! vdd! 366 361 353 357 PG_Blk $T=24800 210235 1 270 $X=11790 $Y=198830
X11 A20_b A20 B20 B20_b gnd! vdd! 386 381 373 377 PG_Blk $T=38850 210235 1 270 $X=25840 $Y=198830
X12 A19_b A19 B19 B19_b gnd! vdd! 406 401 393 397 PG_Blk $T=52900 210235 1 270 $X=39890 $Y=198830
X13 A18_b A18 B18 B18_b gnd! vdd! 425 420 412 416 PG_Blk $T=66950 210235 1 270 $X=53940 $Y=198830
X14 A17_b A17 B17 B17_b gnd! vdd! 446 441 433 437 PG_Blk $T=81000 210235 1 270 $X=67990 $Y=198830
X15 A16_b A16 B16 B16_b gnd! vdd! 466 461 453 457 PG_Blk $T=95050 210235 1 270 $X=82040 $Y=198830
X16 A15_b A15 B15 B15_b gnd! vdd! 484 479 471 475 PG_Blk $T=109100 210235 1 270 $X=96090 $Y=198830
X17 A14_b A14 B14 B14_b gnd! vdd! 497 494 488 491 PG_Blk $T=123150 210235 1 270 $X=110140 $Y=198830
X18 A13_b A13 B13 B13_b gnd! vdd! 509 506 500 503 PG_Blk $T=137200 210235 1 270 $X=124190 $Y=198830
X19 A12_b A12 B12 B12_b gnd! vdd! 521 518 512 515 PG_Blk $T=151250 210235 1 270 $X=138240 $Y=198830
X20 A11_b A11 B11 B11_b gnd! vdd! 533 530 524 527 PG_Blk $T=165300 210235 1 270 $X=152290 $Y=198830
X21 A10_b A10 B10 B10_b gnd! vdd! 545 542 536 539 PG_Blk $T=179350 210235 1 270 $X=166340 $Y=198830
X22 A9_b A9 B9 B9_b gnd! vdd! 557 554 548 551 PG_Blk $T=193400 210235 1 270 $X=180390 $Y=198830
X23 A8_b A8 B8 B8_b gnd! vdd! 569 566 560 563 PG_Blk $T=207450 210235 1 270 $X=194440 $Y=198830
X24 A7_b A7 B7 B7_b gnd! vdd! 581 578 572 575 PG_Blk $T=221500 210235 1 270 $X=208490 $Y=198830
X25 A6_b A6 B6 B6_b gnd! vdd! 589 587 583 585 PG_Blk $T=235550 210235 1 270 $X=222540 $Y=198830
X26 A5_b A5 B5 B5_b gnd! vdd! 597 595 591 593 PG_Blk $T=249600 210235 1 270 $X=236590 $Y=198830
X27 A4_b A4 B4 B4_b gnd! vdd! 605 603 599 601 PG_Blk $T=263650 210235 1 270 $X=250640 $Y=198830
X28 A3_b A3 B3 B3_b gnd! vdd! 613 611 607 609 PG_Blk $T=277700 210235 1 270 $X=264690 $Y=198830
X29 A2_b A2 B2 B2_b gnd! vdd! 617 616 614 615 PG_Blk $T=291750 210235 1 270 $X=278740 $Y=198830
X30 A1_b A1 B1 B1_b gnd! vdd! 621 620 618 619 PG_Blk $T=305800 210235 1 270 $X=292790 $Y=198830
X31 A0_b A0 B0 B0_b gnd! vdd! 485 480 745 622 PG_Blk $T=319850 210235 1 270 $X=306840 $Y=198830
X32 S31 167 168 169 166 gnd! vdd! SP_XOR $T=-128585 36780 1 270 $X=-132190 $Y=30380
X33 S30 177 188 189 173 gnd! vdd! SP_XOR $T=-114580 36780 1 270 $X=-118185 $Y=30380
X34 S29 197 208 209 193 gnd! vdd! SP_XOR $T=-100530 36780 1 270 $X=-104135 $Y=30380
X35 S28 217 228 229 213 gnd! vdd! SP_XOR $T=-86480 36780 1 270 $X=-90085 $Y=30380
X36 S27 237 248 249 233 gnd! vdd! SP_XOR $T=-72430 36780 1 270 $X=-76035 $Y=30380
X37 S26 256 268 269 252 gnd! vdd! SP_XOR $T=-58380 36780 1 270 $X=-61985 $Y=30380
X38 S25 277 288 289 273 gnd! vdd! SP_XOR $T=-44330 36780 1 270 $X=-47935 $Y=30380
X39 S24 297 308 309 293 gnd! vdd! SP_XOR $T=-30280 36780 1 270 $X=-33885 $Y=30380
X40 S23 317 328 329 313 gnd! vdd! SP_XOR $T=-16230 36780 1 270 $X=-19835 $Y=30380
X41 S22 336 348 349 332 gnd! vdd! SP_XOR $T=-2180 36780 1 270 $X=-5785 $Y=30380
X42 S21 357 368 369 353 gnd! vdd! SP_XOR $T=11870 36780 1 270 $X=8265 $Y=30380
X43 S20 377 388 389 373 gnd! vdd! SP_XOR $T=25920 36780 1 270 $X=22315 $Y=30380
X44 S19 397 408 409 393 gnd! vdd! SP_XOR $T=39970 36780 1 270 $X=36365 $Y=30380
X45 S18 416 428 429 412 gnd! vdd! SP_XOR $T=54020 36780 1 270 $X=50415 $Y=30380
X46 S17 437 448 449 433 gnd! vdd! SP_XOR $T=68070 36780 1 270 $X=64465 $Y=30380
X47 S16 457 182 187 453 gnd! vdd! SP_XOR $T=82120 36780 1 270 $X=78515 $Y=30380
X48 S15 475 202 207 471 gnd! vdd! SP_XOR $T=96170 36780 1 270 $X=92565 $Y=30380
X49 S14 491 222 227 488 gnd! vdd! SP_XOR $T=110220 36780 1 270 $X=106615 $Y=30380
X50 S13 503 242 247 500 gnd! vdd! SP_XOR $T=124270 36780 1 270 $X=120665 $Y=30380
X51 S12 515 262 267 512 gnd! vdd! SP_XOR $T=138320 36780 1 270 $X=134715 $Y=30380
X52 S11 527 282 287 524 gnd! vdd! SP_XOR $T=152370 36780 1 270 $X=148765 $Y=30380
X53 S10 539 302 307 536 gnd! vdd! SP_XOR $T=166420 36780 1 270 $X=162815 $Y=30380
X54 S9 551 322 327 548 gnd! vdd! SP_XOR $T=180470 36780 1 270 $X=176865 $Y=30380
X55 S8 563 342 347 560 gnd! vdd! SP_XOR $T=194520 36780 1 270 $X=190915 $Y=30380
X56 S7 575 362 367 572 gnd! vdd! SP_XOR $T=208570 36780 1 270 $X=204965 $Y=30380
X57 S6 585 382 387 583 gnd! vdd! SP_XOR $T=222620 36780 1 270 $X=219015 $Y=30380
X58 S5 593 402 407 591 gnd! vdd! SP_XOR $T=236670 36780 1 270 $X=233065 $Y=30380
X59 S4 601 422 427 599 gnd! vdd! SP_XOR $T=250720 36780 1 270 $X=247115 $Y=30380
X60 S3 609 442 447 607 gnd! vdd! SP_XOR $T=264770 36780 1 270 $X=261165 $Y=30380
X61 S2 615 462 467 614 gnd! vdd! SP_XOR $T=278820 36780 1 270 $X=275215 $Y=30380
X62 S1 619 480 485 618 gnd! vdd! SP_XOR $T=295545 36780 1 270 $X=291940 $Y=30380
X63 S0 622 GND_PC VDD_PC 745 gnd! vdd! SP_XOR $T=309595 36780 1 270 $X=305990 $Y=30380
X64 187 182 636 635 634 633 gnd! OV gnd! vdd! GREY_CELL $T=-119165 54165 1 270 $X=-123535 $Y=45830
X65 207 202 653 652 651 650 169 168 gnd! vdd! GREY_CELL $T=-105115 54165 1 270 $X=-109485 $Y=45830
X66 227 222 666 665 664 663 189 188 gnd! vdd! GREY_CELL $T=-91065 54165 1 270 $X=-95435 $Y=45830
X67 247 242 678 677 676 675 209 208 gnd! vdd! GREY_CELL $T=-77015 54165 1 270 $X=-81385 $Y=45830
X68 267 262 687 686 685 684 229 228 gnd! vdd! GREY_CELL $T=-62965 54165 1 270 $X=-67335 $Y=45830
X69 287 282 695 694 693 692 249 248 gnd! vdd! GREY_CELL $T=-48915 54165 1 270 $X=-53285 $Y=45830
X70 307 302 703 702 701 700 269 268 gnd! vdd! GREY_CELL $T=-34865 54165 1 270 $X=-39235 $Y=45830
X71 327 322 711 710 709 708 289 288 gnd! vdd! GREY_CELL $T=-20815 54165 1 270 $X=-25185 $Y=45830
X72 347 342 716 715 714 713 309 308 gnd! vdd! GREY_CELL $T=-6765 54165 1 270 $X=-11135 $Y=45830
X73 367 362 720 719 718 717 329 328 gnd! vdd! GREY_CELL $T=7285 54165 1 270 $X=2915 $Y=45830
X74 387 382 724 723 722 721 349 348 gnd! vdd! GREY_CELL $T=21335 54165 1 270 $X=16965 $Y=45830
X75 407 402 728 727 726 725 369 368 gnd! vdd! GREY_CELL $T=35385 54165 1 270 $X=31015 $Y=45830
X76 427 422 732 731 730 729 389 388 gnd! vdd! GREY_CELL $T=49435 54165 1 270 $X=45065 $Y=45830
X77 447 442 736 735 734 733 409 408 gnd! vdd! GREY_CELL $T=63485 54165 1 270 $X=59115 $Y=45830
X78 467 462 740 739 738 737 429 428 gnd! vdd! GREY_CELL $T=77535 54165 1 270 $X=73165 $Y=45830
X79 485 480 744 743 742 741 449 448 gnd! vdd! GREY_CELL $T=91585 54165 1 270 $X=87215 $Y=45830
X80 347 342 343 338 334 330 187 182 gnd! vdd! GREY_CELL $T=105635 95560 1 270 $X=101265 $Y=87225
X81 367 362 363 358 354 350 207 202 gnd! vdd! GREY_CELL $T=119685 95560 1 270 $X=115315 $Y=87225
X82 387 382 383 378 374 370 227 222 gnd! vdd! GREY_CELL $T=133735 95560 1 270 $X=129365 $Y=87225
X83 407 402 403 398 394 390 247 242 gnd! vdd! GREY_CELL $T=147785 95560 1 270 $X=143415 $Y=87225
X84 427 422 423 418 414 410 267 262 gnd! vdd! GREY_CELL $T=161835 95560 1 270 $X=157465 $Y=87225
X85 447 442 443 438 434 430 287 282 gnd! vdd! GREY_CELL $T=175885 95560 1 270 $X=171515 $Y=87225
X86 467 462 463 458 454 450 307 302 gnd! vdd! GREY_CELL $T=189935 95560 1 270 $X=185565 $Y=87225
X87 485 480 481 476 472 468 327 322 gnd! vdd! GREY_CELL $T=203985 95560 1 270 $X=199615 $Y=87225
X88 427 422 543 540 537 534 347 342 gnd! vdd! GREY_CELL $T=218035 137105 1 270 $X=213665 $Y=128770
X89 447 442 555 552 549 546 367 362 gnd! vdd! GREY_CELL $T=232085 137105 1 270 $X=227715 $Y=128770
X90 467 462 567 564 561 558 387 382 gnd! vdd! GREY_CELL $T=246135 137105 1 270 $X=241765 $Y=128770
X91 485 480 579 576 573 570 407 402 gnd! vdd! GREY_CELL $T=260185 137105 1 270 $X=255815 $Y=128770
X92 467 462 604 602 600 598 427 422 gnd! vdd! GREY_CELL $T=274235 169410 1 270 $X=269865 $Y=161075
X93 485 480 612 610 608 606 447 442 gnd! vdd! GREY_CELL $T=288285 169410 1 270 $X=283915 $Y=161075
X94 485 480 621 620 619 618 467 462 gnd! vdd! GREY_CELL $T=302445 192410 1 270 $X=298075 $Y=184075
X95 170 174 629 637 623 626 183 gnd! vdd! 178 636 635 634 633 BLACK_CELL $T=-113550 93125 1 270 $X=-128595 $Y=84525
X96 171 175 630 638 624 627 184 gnd! vdd! 179 637 629 626 623 BLACK_CELL $T=-113550 134670 1 270 $X=-128595 $Y=126070
X97 172 176 631 639 625 628 185 gnd! vdd! 180 638 630 627 624 BLACK_CELL $T=-113550 166970 1 270 $X=-128595 $Y=158370
X98 173 177 632 640 166 167 186 gnd! vdd! 181 639 631 628 625 BLACK_CELL $T=-113550 189975 1 270 $X=-128595 $Y=181375
X99 190 194 647 654 641 644 203 gnd! vdd! 198 653 652 651 650 BLACK_CELL $T=-99500 93125 1 270 $X=-114545 $Y=84525
X100 191 195 648 655 642 645 204 gnd! vdd! 199 654 647 644 641 BLACK_CELL $T=-99500 134670 1 270 $X=-114545 $Y=126070
X101 192 196 649 656 643 646 205 gnd! vdd! 200 655 648 645 642 BLACK_CELL $T=-99500 166970 1 270 $X=-114545 $Y=158370
X102 193 197 181 186 173 177 206 gnd! vdd! 201 656 649 646 643 BLACK_CELL $T=-99500 189975 1 270 $X=-114545 $Y=181375
X103 210 214 661 667 657 659 223 gnd! vdd! 218 666 665 664 663 BLACK_CELL $T=-85450 93125 1 270 $X=-100495 $Y=84525
X104 211 215 662 668 658 660 224 gnd! vdd! 219 667 661 659 657 BLACK_CELL $T=-85450 134670 1 270 $X=-100495 $Y=126070
X105 212 216 180 185 172 176 225 gnd! vdd! 220 668 662 660 658 BLACK_CELL $T=-85450 166970 1 270 $X=-100495 $Y=158370
X106 213 217 201 206 193 197 226 gnd! vdd! 221 185 180 176 172 BLACK_CELL $T=-85450 189975 1 270 $X=-100495 $Y=181375
X107 230 234 673 679 669 671 243 gnd! vdd! 238 678 677 676 675 BLACK_CELL $T=-71400 93125 1 270 $X=-86445 $Y=84525
X108 231 235 674 680 670 672 244 gnd! vdd! 239 679 673 671 669 BLACK_CELL $T=-71400 134670 1 270 $X=-86445 $Y=126070
X109 232 236 200 205 192 196 245 gnd! vdd! 240 680 674 672 670 BLACK_CELL $T=-71400 166970 1 270 $X=-86445 $Y=158370
X110 233 237 221 226 213 217 246 gnd! vdd! 241 205 200 196 192 BLACK_CELL $T=-71400 189975 1 270 $X=-86445 $Y=181375
X111 250 254 683 688 681 682 263 gnd! vdd! 258 687 686 685 684 BLACK_CELL $T=-57350 93125 1 270 $X=-72395 $Y=84525
X112 251 255 179 184 171 175 264 gnd! vdd! 259 688 683 682 681 BLACK_CELL $T=-57350 134670 1 270 $X=-72395 $Y=126070
X113 253 257 220 225 212 216 266 gnd! vdd! 261 184 179 175 171 BLACK_CELL $T=-57350 166970 1 270 $X=-72395 $Y=158370
X114 252 256 241 246 233 237 265 gnd! vdd! 260 225 220 216 212 BLACK_CELL $T=-57350 189975 1 270 $X=-72395 $Y=181375
X115 270 274 691 696 689 690 283 gnd! vdd! 278 695 694 693 692 BLACK_CELL $T=-43300 93125 1 270 $X=-58345 $Y=84525
X116 271 275 199 204 191 195 284 gnd! vdd! 279 696 691 690 689 BLACK_CELL $T=-43300 134670 1 270 $X=-58345 $Y=126070
X117 272 276 240 245 232 236 285 gnd! vdd! 280 204 199 195 191 BLACK_CELL $T=-43300 166970 1 270 $X=-58345 $Y=158370
X118 273 277 260 265 252 256 286 gnd! vdd! 281 245 240 236 232 BLACK_CELL $T=-43300 189975 1 270 $X=-58345 $Y=181375
X119 290 294 699 704 697 698 303 gnd! vdd! 298 703 702 701 700 BLACK_CELL $T=-29250 93125 1 270 $X=-44295 $Y=84525
X120 291 295 219 224 211 215 304 gnd! vdd! 299 704 699 698 697 BLACK_CELL $T=-29250 134670 1 270 $X=-44295 $Y=126070
X121 292 296 261 266 253 257 305 gnd! vdd! 300 224 219 215 211 BLACK_CELL $T=-29250 166970 1 270 $X=-44295 $Y=158370
X122 293 297 281 286 273 277 306 gnd! vdd! 301 266 261 257 253 BLACK_CELL $T=-29250 189975 1 270 $X=-44295 $Y=181375
X123 310 314 707 712 705 706 323 gnd! vdd! 318 711 710 709 708 BLACK_CELL $T=-15200 93125 1 270 $X=-30245 $Y=84525
X124 311 315 239 244 231 235 324 gnd! vdd! 319 712 707 706 705 BLACK_CELL $T=-15200 134670 1 270 $X=-30245 $Y=126070
X125 312 316 280 285 272 276 325 gnd! vdd! 320 244 239 235 231 BLACK_CELL $T=-15200 166970 1 270 $X=-30245 $Y=158370
X126 313 317 301 306 293 297 326 gnd! vdd! 321 285 280 276 272 BLACK_CELL $T=-15200 189975 1 270 $X=-30245 $Y=181375
X127 330 334 178 183 170 174 343 gnd! vdd! 338 716 715 714 713 BLACK_CELL $T=-1150 93125 1 270 $X=-16195 $Y=84525
X128 331 335 259 264 251 255 344 gnd! vdd! 339 183 178 174 170 BLACK_CELL $T=-1150 134670 1 270 $X=-16195 $Y=126070
X129 333 337 300 305 292 296 346 gnd! vdd! 341 264 259 255 251 BLACK_CELL $T=-1150 166970 1 270 $X=-16195 $Y=158370
X130 332 336 321 326 313 317 345 gnd! vdd! 340 305 300 296 292 BLACK_CELL $T=-1150 189975 1 270 $X=-16195 $Y=181375
X131 350 354 198 203 190 194 363 gnd! vdd! 358 720 719 718 717 BLACK_CELL $T=12900 93125 1 270 $X=-2145 $Y=84525
X132 351 355 279 284 271 275 364 gnd! vdd! 359 203 198 194 190 BLACK_CELL $T=12900 134670 1 270 $X=-2145 $Y=126070
X133 352 356 320 325 312 316 365 gnd! vdd! 360 284 279 275 271 BLACK_CELL $T=12900 166970 1 270 $X=-2145 $Y=158370
X134 353 357 340 345 332 336 366 gnd! vdd! 361 325 320 316 312 BLACK_CELL $T=12900 189975 1 270 $X=-2145 $Y=181375
X135 370 374 218 223 210 214 383 gnd! vdd! 378 724 723 722 721 BLACK_CELL $T=26950 93125 1 270 $X=11905 $Y=84525
X136 371 375 299 304 291 295 384 gnd! vdd! 379 223 218 214 210 BLACK_CELL $T=26950 134670 1 270 $X=11905 $Y=126070
X137 372 376 341 346 333 337 385 gnd! vdd! 380 304 299 295 291 BLACK_CELL $T=26950 166970 1 270 $X=11905 $Y=158370
X138 373 377 361 366 353 357 386 gnd! vdd! 381 346 341 337 333 BLACK_CELL $T=26950 189975 1 270 $X=11905 $Y=181375
X139 390 394 238 243 230 234 403 gnd! vdd! 398 728 727 726 725 BLACK_CELL $T=41000 93125 1 270 $X=25955 $Y=84525
X140 391 395 319 324 311 315 404 gnd! vdd! 399 243 238 234 230 BLACK_CELL $T=41000 134670 1 270 $X=25955 $Y=126070
X141 392 396 360 365 352 356 405 gnd! vdd! 400 324 319 315 311 BLACK_CELL $T=41000 166970 1 270 $X=25955 $Y=158370
X142 393 397 381 386 373 377 406 gnd! vdd! 401 365 360 356 352 BLACK_CELL $T=41000 189975 1 270 $X=25955 $Y=181375
X143 410 414 258 263 250 254 423 gnd! vdd! 418 732 731 730 729 BLACK_CELL $T=55050 93125 1 270 $X=40005 $Y=84525
X144 411 415 339 344 331 335 424 gnd! vdd! 419 263 258 254 250 BLACK_CELL $T=55050 134670 1 270 $X=40005 $Y=126070
X145 413 417 380 385 372 376 426 gnd! vdd! 421 344 339 335 331 BLACK_CELL $T=55050 166970 1 270 $X=40005 $Y=158370
X146 412 416 401 406 393 397 425 gnd! vdd! 420 385 380 376 372 BLACK_CELL $T=55050 189975 1 270 $X=40005 $Y=181375
X147 430 434 278 283 270 274 443 gnd! vdd! 438 736 735 734 733 BLACK_CELL $T=69100 93125 1 270 $X=54055 $Y=84525
X148 431 435 359 364 351 355 444 gnd! vdd! 439 283 278 274 270 BLACK_CELL $T=69100 134670 1 270 $X=54055 $Y=126070
X149 432 436 400 405 392 396 445 gnd! vdd! 440 364 359 355 351 BLACK_CELL $T=69100 166970 1 270 $X=54055 $Y=158370
X150 433 437 420 425 412 416 446 gnd! vdd! 441 405 400 396 392 BLACK_CELL $T=69100 189975 1 270 $X=54055 $Y=181375
X151 450 454 298 303 290 294 463 gnd! vdd! 458 740 739 738 737 BLACK_CELL $T=83150 93125 1 270 $X=68105 $Y=84525
X152 451 455 379 384 371 375 464 gnd! vdd! 459 303 298 294 290 BLACK_CELL $T=83150 134670 1 270 $X=68105 $Y=126070
X153 452 456 421 426 413 417 465 gnd! vdd! 460 384 379 375 371 BLACK_CELL $T=83150 166970 1 270 $X=68105 $Y=158370
X154 453 457 441 446 433 437 466 gnd! vdd! 461 426 421 417 413 BLACK_CELL $T=83150 189975 1 270 $X=68105 $Y=181375
X155 468 472 318 323 310 314 481 gnd! vdd! 476 744 743 742 741 BLACK_CELL $T=97200 93125 1 270 $X=82155 $Y=84525
X156 469 473 399 404 391 395 482 gnd! vdd! 477 323 318 314 310 BLACK_CELL $T=97200 134670 1 270 $X=82155 $Y=126070
X157 470 474 440 445 432 436 483 gnd! vdd! 478 404 399 395 391 BLACK_CELL $T=97200 166970 1 270 $X=82155 $Y=158370
X158 471 475 461 466 453 457 484 gnd! vdd! 479 445 440 436 432 BLACK_CELL $T=97200 189975 1 270 $X=82155 $Y=181375
X159 486 489 419 424 411 415 495 gnd! vdd! 492 343 338 334 330 BLACK_CELL $T=111250 134670 1 270 $X=96205 $Y=126070
X160 487 490 460 465 452 456 496 gnd! vdd! 493 424 419 415 411 BLACK_CELL $T=111250 166970 1 270 $X=96205 $Y=158370
X161 488 491 479 484 471 475 497 gnd! vdd! 494 465 460 456 452 BLACK_CELL $T=111250 189975 1 270 $X=96205 $Y=181375
X162 498 501 439 444 431 435 507 gnd! vdd! 504 363 358 354 350 BLACK_CELL $T=125300 134670 1 270 $X=110255 $Y=126070
X163 499 502 478 483 470 474 508 gnd! vdd! 505 444 439 435 431 BLACK_CELL $T=125300 166970 1 270 $X=110255 $Y=158370
X164 500 503 494 497 488 491 509 gnd! vdd! 506 483 478 474 470 BLACK_CELL $T=125300 189975 1 270 $X=110255 $Y=181375
X165 510 513 459 464 451 455 519 gnd! vdd! 516 383 378 374 370 BLACK_CELL $T=139350 134670 1 270 $X=124305 $Y=126070
X166 511 514 493 496 487 490 520 gnd! vdd! 517 464 459 455 451 BLACK_CELL $T=139350 166970 1 270 $X=124305 $Y=158370
X167 512 515 506 509 500 503 521 gnd! vdd! 518 496 493 490 487 BLACK_CELL $T=139350 189975 1 270 $X=124305 $Y=181375
X168 522 525 477 482 469 473 531 gnd! vdd! 528 403 398 394 390 BLACK_CELL $T=153400 134670 1 270 $X=138355 $Y=126070
X169 523 526 505 508 499 502 532 gnd! vdd! 529 482 477 473 469 BLACK_CELL $T=153400 166970 1 270 $X=138355 $Y=158370
X170 524 527 518 521 512 515 533 gnd! vdd! 530 508 505 502 499 BLACK_CELL $T=153400 189975 1 270 $X=138355 $Y=181375
X171 534 537 492 495 486 489 543 gnd! vdd! 540 423 418 414 410 BLACK_CELL $T=167450 134670 1 270 $X=152405 $Y=126070
X172 535 538 517 520 511 514 544 gnd! vdd! 541 495 492 489 486 BLACK_CELL $T=167450 166970 1 270 $X=152405 $Y=158370
X173 536 539 530 533 524 527 545 gnd! vdd! 542 520 517 514 511 BLACK_CELL $T=167450 189975 1 270 $X=152405 $Y=181375
X174 546 549 504 507 498 501 555 gnd! vdd! 552 443 438 434 430 BLACK_CELL $T=181500 134670 1 270 $X=166455 $Y=126070
X175 547 550 529 532 523 526 556 gnd! vdd! 553 507 504 501 498 BLACK_CELL $T=181500 166970 1 270 $X=166455 $Y=158370
X176 548 551 542 545 536 539 557 gnd! vdd! 554 532 529 526 523 BLACK_CELL $T=181500 189975 1 270 $X=166455 $Y=181375
X177 558 561 516 519 510 513 567 gnd! vdd! 564 463 458 454 450 BLACK_CELL $T=195550 134670 1 270 $X=180505 $Y=126070
X178 559 562 541 544 535 538 568 gnd! vdd! 565 519 516 513 510 BLACK_CELL $T=195550 166970 1 270 $X=180505 $Y=158370
X179 560 563 554 557 548 551 569 gnd! vdd! 566 544 541 538 535 BLACK_CELL $T=195550 189975 1 270 $X=180505 $Y=181375
X180 570 573 528 531 522 525 579 gnd! vdd! 576 481 476 472 468 BLACK_CELL $T=209600 134670 1 270 $X=194555 $Y=126070
X181 571 574 553 556 547 550 580 gnd! vdd! 577 531 528 525 522 BLACK_CELL $T=209600 166970 1 270 $X=194555 $Y=158370
X182 572 575 566 569 560 563 581 gnd! vdd! 578 556 553 550 547 BLACK_CELL $T=209600 189975 1 270 $X=194555 $Y=181375
X183 582 584 565 568 559 562 588 gnd! vdd! 586 543 540 537 534 BLACK_CELL $T=223650 166970 1 270 $X=208605 $Y=158370
X184 583 585 578 581 572 575 589 gnd! vdd! 587 568 565 562 559 BLACK_CELL $T=223650 189975 1 270 $X=208605 $Y=181375
X185 590 592 577 580 571 574 596 gnd! vdd! 594 555 552 549 546 BLACK_CELL $T=237700 166970 1 270 $X=222655 $Y=158370
X186 591 593 587 589 583 585 597 gnd! vdd! 595 580 577 574 571 BLACK_CELL $T=237700 189975 1 270 $X=222655 $Y=181375
X187 598 600 586 588 582 584 604 gnd! vdd! 602 567 564 561 558 BLACK_CELL $T=251750 166970 1 270 $X=236705 $Y=158370
X188 599 601 595 597 591 593 605 gnd! vdd! 603 588 586 584 582 BLACK_CELL $T=251750 189975 1 270 $X=236705 $Y=181375
X189 606 608 594 596 590 592 612 gnd! vdd! 610 579 576 573 570 BLACK_CELL $T=265800 166970 1 270 $X=250755 $Y=158370
X190 607 609 603 605 599 601 613 gnd! vdd! 611 596 594 592 590 BLACK_CELL $T=265800 189975 1 270 $X=250755 $Y=181375
X191 614 615 611 613 607 609 617 gnd! vdd! 616 604 602 600 598 BLACK_CELL $T=279850 189975 1 270 $X=264805 $Y=181375
X192 618 619 616 617 614 615 621 gnd! vdd! 620 612 610 608 606 BLACK_CELL $T=293900 189975 1 270 $X=278855 $Y=181375
.ENDS
***************************************
.SUBCKT SP_42CSA_DR gnd! vdd! Z31 Z31_b C31 C31_b Z30 Z30_b C30 C30_b Z29 Z29_b C29 C29_b Z28 Z28_b C28 C28_b Z27 Z27_b
+ C27 C27_b Z26 Z26_b C26 C26_b Z25 Z25_b C25 C25_b Z24 Z24_b C24 C24_b Z23 Z23_b C23 C23_b Z22 Z22_b
+ C22 C22_b Z21 Z21_b C21 C21_b Z20 Z20_b C20 C20_b Z19 Z19_b C19 C19_b Z18 Z18_b C18 C18_b Z17 Z17_b
+ C17 C17_b Z16 Z16_b C16 C16_b Z15 Z15_b C15 C15_b Z14 Z14_b C14 C14_b Z13 Z13_b C13 C13_b Z12 Z12_b
+ C12 C12_b Z11 Z11_b C11 C11_b Z10 Z10_b C10 C10_b Z9 Z9_b C9 C9_b Z8 Z8_b C8 C8_b Z7 Z7_b
+ C7 C7_b Z6 Z6_b C6 C6_b Z5 Z5_b C5 C5_b Z4 Z4_b C4 C4_b Z3 Z3_b C3 C3_b Z2 Z2_b
+ C2 C2_b Z1 Z1_b C1 C1_b Z0 Z0_b W31 W31_b X31 X31_b Y31 Y31_b S31 S31_b W30 W30_b X30 X30_b
+ Y30 Y30_b S30 S30_b W29 W29_b X29 X29_b Y29 Y29_b S29 S29_b W28 W28_b X28 X28_b Y28 Y28_b S28 S28_b
+ W27 W27_b X27 X27_b Y27 Y27_b S27 S27_b W26 W26_b X26 X26_b Y26 Y26_b S26 S26_b W25 W25_b X25 X25_b
+ Y25 Y25_b S25 S25_b W24 W24_b X24 X24_b Y24 Y24_b S24 S24_b W23 W23_b X23 X23_b Y23 Y23_b S23 S23_b
+ W22 W22_b X22 X22_b Y22 Y22_b S22 S22_b W21 W21_b X21 X21_b Y21 Y21_b S21 S21_b W20 W20_b X20 X20_b
+ Y20 Y20_b S20 S20_b W19 W19_b X19 X19_b Y19 Y19_b S19 S19_b W18 W18_b X18 X18_b Y18 Y18_b S18 S18_b
+ W17 W17_b X17 X17_b Y17 Y17_b S17 S17_b W16 W16_b X16 X16_b Y16 Y16_b S16 S16_b W15 W15_b X15 X15_b
+ Y15 Y15_b S15 S15_b W14 W14_b X14 X14_b Y14 Y14_b S14 S14_b W13 W13_b X13 X13_b Y13 Y13_b S13 S13_b
+ W12 W12_b X12 X12_b Y12 Y12_b S12 S12_b W11 W11_b X11 X11_b Y11 Y11_b S11 S11_b W10 W10_b X10 X10_b
+ Y10 Y10_b S10 S10_b W9 W9_b X9 X9_b Y9 Y9_b S9 S9_b W8 W8_b X8 X8_b Y8 Y8_b S8 S8_b
+ W7 W7_b X7 X7_b Y7 Y7_b S7 S7_b W6 W6_b X6 X6_b Y6 Y6_b S6 S6_b W5 W5_b X5 X5_b
+ Y5 Y5_b S5 S5_b W4 W4_b X4 X4_b Y4 Y4_b S4 S4_b W3 W3_b X3 X3_b Y3 Y3_b S3 S3_b
+ W2 W2_b X2 X2_b Y2 Y2_b S2 S2_b W1 W1_b X1 X1_b Y1 Y1_b S1 S1_b W0 W0_b X0 X0_b
+ Y0 Y0_b S0 S0_b
** N=510 EP=384 IP=830 FDC=3456
X62 vdd! 198 Z31 5 200 gnd! Z31_b 6 S31 S31_b gnd! gnd! SP_FA_DR $T=-107445 128150 0 0 $X=-103125 $Y=128650
X63 vdd! W31 X31 Y31 W31_b gnd! X31_b Y31_b 198 200 gnd! gnd! SP_FA_DR $T=-107445 148705 0 0 $X=-103125 $Y=149205
X64 vdd! 208 Z30 11 210 gnd! Z30_b 12 S30 S30_b C31 C31_b SP_FA_DR $T=-89485 128150 0 0 $X=-85165 $Y=128650
X65 vdd! W30 X30 Y30 W30_b gnd! X30_b Y30_b 208 210 5 6 SP_FA_DR $T=-89485 148705 0 0 $X=-85165 $Y=149205
X66 vdd! 218 Z29 17 220 gnd! Z29_b 18 S29 S29_b C30 C30_b SP_FA_DR $T=-71525 128150 0 0 $X=-67205 $Y=128650
X67 vdd! W29 X29 Y29 W29_b gnd! X29_b Y29_b 218 220 11 12 SP_FA_DR $T=-71525 148705 0 0 $X=-67205 $Y=149205
X68 vdd! 228 Z28 23 230 gnd! Z28_b 24 S28 S28_b C29 C29_b SP_FA_DR $T=-53565 128150 0 0 $X=-49245 $Y=128650
X69 vdd! W28 X28 Y28 W28_b gnd! X28_b Y28_b 228 230 17 18 SP_FA_DR $T=-53565 148705 0 0 $X=-49245 $Y=149205
X70 vdd! 238 Z27 29 240 gnd! Z27_b 30 S27 S27_b C28 C28_b SP_FA_DR $T=-35605 128150 0 0 $X=-31285 $Y=128650
X71 vdd! W27 X27 Y27 W27_b gnd! X27_b Y27_b 238 240 23 24 SP_FA_DR $T=-35605 148705 0 0 $X=-31285 $Y=149205
X72 vdd! 248 Z26 35 250 gnd! Z26_b 36 S26 S26_b C27 C27_b SP_FA_DR $T=-17645 128150 0 0 $X=-13325 $Y=128650
X73 vdd! W26 X26 Y26 W26_b gnd! X26_b Y26_b 248 250 29 30 SP_FA_DR $T=-17645 148705 0 0 $X=-13325 $Y=149205
X74 vdd! 258 Z25 41 260 gnd! Z25_b 42 S25 S25_b C26 C26_b SP_FA_DR $T=315 128150 0 0 $X=4635 $Y=128650
X75 vdd! W25 X25 Y25 W25_b gnd! X25_b Y25_b 258 260 35 36 SP_FA_DR $T=315 148705 0 0 $X=4635 $Y=149205
X76 vdd! 268 Z24 47 270 gnd! Z24_b 48 S24 S24_b C25 C25_b SP_FA_DR $T=18275 128150 0 0 $X=22595 $Y=128650
X77 vdd! W24 X24 Y24 W24_b gnd! X24_b Y24_b 268 270 41 42 SP_FA_DR $T=18275 148705 0 0 $X=22595 $Y=149205
X78 vdd! 278 Z23 53 280 gnd! Z23_b 54 S23 S23_b C24 C24_b SP_FA_DR $T=36235 128150 0 0 $X=40555 $Y=128650
X79 vdd! W23 X23 Y23 W23_b gnd! X23_b Y23_b 278 280 47 48 SP_FA_DR $T=36235 148705 0 0 $X=40555 $Y=149205
X80 vdd! 288 Z22 59 290 gnd! Z22_b 60 S22 S22_b C23 C23_b SP_FA_DR $T=54195 128150 0 0 $X=58515 $Y=128650
X81 vdd! W22 X22 Y22 W22_b gnd! X22_b Y22_b 288 290 53 54 SP_FA_DR $T=54195 148705 0 0 $X=58515 $Y=149205
X82 vdd! 298 Z21 65 300 gnd! Z21_b 66 S21 S21_b C22 C22_b SP_FA_DR $T=72155 128150 0 0 $X=76475 $Y=128650
X83 vdd! W21 X21 Y21 W21_b gnd! X21_b Y21_b 298 300 59 60 SP_FA_DR $T=72155 148705 0 0 $X=76475 $Y=149205
X84 vdd! 308 Z20 71 310 gnd! Z20_b 72 S20 S20_b C21 C21_b SP_FA_DR $T=90115 128150 0 0 $X=94435 $Y=128650
X85 vdd! W20 X20 Y20 W20_b gnd! X20_b Y20_b 308 310 65 66 SP_FA_DR $T=90115 148705 0 0 $X=94435 $Y=149205
X86 vdd! 318 Z19 77 320 gnd! Z19_b 78 S19 S19_b C20 C20_b SP_FA_DR $T=108075 128150 0 0 $X=112395 $Y=128650
X87 vdd! W19 X19 Y19 W19_b gnd! X19_b Y19_b 318 320 71 72 SP_FA_DR $T=108075 148705 0 0 $X=112395 $Y=149205
X88 vdd! 328 Z18 83 330 gnd! Z18_b 84 S18 S18_b C19 C19_b SP_FA_DR $T=126035 128150 0 0 $X=130355 $Y=128650
X89 vdd! W18 X18 Y18 W18_b gnd! X18_b Y18_b 328 330 77 78 SP_FA_DR $T=126035 148705 0 0 $X=130355 $Y=149205
X90 vdd! 338 Z17 89 340 gnd! Z17_b 90 S17 S17_b C18 C18_b SP_FA_DR $T=143995 128150 0 0 $X=148315 $Y=128650
X91 vdd! W17 X17 Y17 W17_b gnd! X17_b Y17_b 338 340 83 84 SP_FA_DR $T=143995 148705 0 0 $X=148315 $Y=149205
X92 vdd! 348 Z16 95 350 gnd! Z16_b 96 S16 S16_b C17 C17_b SP_FA_DR $T=161955 128150 0 0 $X=166275 $Y=128650
X93 vdd! W16 X16 Y16 W16_b gnd! X16_b Y16_b 348 350 89 90 SP_FA_DR $T=161955 148705 0 0 $X=166275 $Y=149205
X94 vdd! 358 Z15 101 360 gnd! Z15_b 102 S15 S15_b C16 C16_b SP_FA_DR $T=179915 128150 0 0 $X=184235 $Y=128650
X95 vdd! W15 X15 Y15 W15_b gnd! X15_b Y15_b 358 360 95 96 SP_FA_DR $T=179915 148705 0 0 $X=184235 $Y=149205
X96 vdd! 368 Z14 107 370 gnd! Z14_b 108 S14 S14_b C15 C15_b SP_FA_DR $T=197875 128150 0 0 $X=202195 $Y=128650
X97 vdd! W14 X14 Y14 W14_b gnd! X14_b Y14_b 368 370 101 102 SP_FA_DR $T=197875 148705 0 0 $X=202195 $Y=149205
X98 vdd! 378 Z13 113 380 gnd! Z13_b 114 S13 S13_b C14 C14_b SP_FA_DR $T=215835 128150 0 0 $X=220155 $Y=128650
X99 vdd! W13 X13 Y13 W13_b gnd! X13_b Y13_b 378 380 107 108 SP_FA_DR $T=215835 148705 0 0 $X=220155 $Y=149205
X100 vdd! 388 Z12 119 390 gnd! Z12_b 120 S12 S12_b C13 C13_b SP_FA_DR $T=233795 128150 0 0 $X=238115 $Y=128650
X101 vdd! W12 X12 Y12 W12_b gnd! X12_b Y12_b 388 390 113 114 SP_FA_DR $T=233795 148705 0 0 $X=238115 $Y=149205
X102 vdd! 398 Z11 125 400 gnd! Z11_b 126 S11 S11_b C12 C12_b SP_FA_DR $T=251755 128150 0 0 $X=256075 $Y=128650
X103 vdd! W11 X11 Y11 W11_b gnd! X11_b Y11_b 398 400 119 120 SP_FA_DR $T=251755 148705 0 0 $X=256075 $Y=149205
X104 vdd! 408 Z10 131 410 gnd! Z10_b 132 S10 S10_b C11 C11_b SP_FA_DR $T=269715 128150 0 0 $X=274035 $Y=128650
X105 vdd! W10 X10 Y10 W10_b gnd! X10_b Y10_b 408 410 125 126 SP_FA_DR $T=269715 148705 0 0 $X=274035 $Y=149205
X106 vdd! 418 Z9 137 420 gnd! Z9_b 138 S9 S9_b C10 C10_b SP_FA_DR $T=287675 128150 0 0 $X=291995 $Y=128650
X107 vdd! W9 X9 Y9 W9_b gnd! X9_b Y9_b 418 420 131 132 SP_FA_DR $T=287675 148705 0 0 $X=291995 $Y=149205
X108 vdd! 428 Z8 143 430 gnd! Z8_b 144 S8 S8_b C9 C9_b SP_FA_DR $T=305635 128150 0 0 $X=309955 $Y=128650
X109 vdd! W8 X8 Y8 W8_b gnd! X8_b Y8_b 428 430 137 138 SP_FA_DR $T=305635 148705 0 0 $X=309955 $Y=149205
X110 vdd! 438 Z7 149 440 gnd! Z7_b 150 S7 S7_b C8 C8_b SP_FA_DR $T=323595 128150 0 0 $X=327915 $Y=128650
X111 vdd! W7 X7 Y7 W7_b gnd! X7_b Y7_b 438 440 143 144 SP_FA_DR $T=323595 148705 0 0 $X=327915 $Y=149205
X112 vdd! 448 Z6 155 450 gnd! Z6_b 156 S6 S6_b C7 C7_b SP_FA_DR $T=341555 128150 0 0 $X=345875 $Y=128650
X113 vdd! W6 X6 Y6 W6_b gnd! X6_b Y6_b 448 450 149 150 SP_FA_DR $T=341555 148705 0 0 $X=345875 $Y=149205
X114 vdd! 458 Z5 161 460 gnd! Z5_b 162 S5 S5_b C6 C6_b SP_FA_DR $T=359515 128150 0 0 $X=363835 $Y=128650
X115 vdd! W5 X5 Y5 W5_b gnd! X5_b Y5_b 458 460 155 156 SP_FA_DR $T=359515 148705 0 0 $X=363835 $Y=149205
X116 vdd! 468 Z4 167 470 gnd! Z4_b 168 S4 S4_b C5 C5_b SP_FA_DR $T=377475 128150 0 0 $X=381795 $Y=128650
X117 vdd! W4 X4 Y4 W4_b gnd! X4_b Y4_b 468 470 161 162 SP_FA_DR $T=377475 148705 0 0 $X=381795 $Y=149205
X118 vdd! 478 Z3 173 480 gnd! Z3_b 174 S3 S3_b C4 C4_b SP_FA_DR $T=395435 128150 0 0 $X=399755 $Y=128650
X119 vdd! W3 X3 Y3 W3_b gnd! X3_b Y3_b 478 480 167 168 SP_FA_DR $T=395435 148705 0 0 $X=399755 $Y=149205
X120 vdd! 488 Z2 179 490 gnd! Z2_b 180 S2 S2_b C3 C3_b SP_FA_DR $T=413395 128150 0 0 $X=417715 $Y=128650
X121 vdd! W2 X2 Y2 W2_b gnd! X2_b Y2_b 488 490 173 174 SP_FA_DR $T=413395 148705 0 0 $X=417715 $Y=149205
X122 vdd! 498 Z1 185 500 gnd! Z1_b 186 S1 S1_b C2 C2_b SP_FA_DR $T=431355 128150 0 0 $X=435675 $Y=128650
X123 vdd! W1 X1 Y1 W1_b gnd! X1_b Y1_b 498 500 179 180 SP_FA_DR $T=431355 148705 0 0 $X=435675 $Y=149205
X124 vdd! 508 Z0 gnd! 510 gnd! Z0_b vdd! S0 S0_b C1 C1_b SP_FA_DR $T=449315 128150 0 0 $X=453635 $Y=128650
X125 vdd! W0 X0 Y0 W0_b gnd! X0_b Y0_b 508 510 185 186 SP_FA_DR $T=449315 148705 0 0 $X=453635 $Y=149205
.ENDS
***************************************
.SUBCKT ICV_5
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT SP_AND3_DR !C !B !A out out_b gnd! vdd! C B A
** N=18 EP=10 IP=4 FDC=22
M0 15 C gnd! gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=5.3325e-14 PD=8.2e-07 PS=9.35e-07 $X=-1085 $Y=-715 $D=1
M1 16 B 15 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=3.78e-14 PD=8.2e-07 PS=8.2e-07 $X=-705 $Y=-715 $D=1
M2 4 A 16 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=4.1175e-14 AS=3.78e-14 PD=8.45e-07 PS=8.2e-07 $X=-325 $Y=-715 $D=1
M3 6 !A gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=900 $Y=-715 $D=1
M4 8 !B gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=2530 $Y=-715 $D=1
M5 14 !C gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=4030 $Y=-715 $D=1
M6 17 6 gnd! gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.835e-14 PD=8.2e-07 PS=7.5e-07 $X=5675 $Y=-935 $D=1
M7 18 8 17 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=3.78e-14 PD=8.2e-07 PS=8.2e-07 $X=6055 $Y=-935 $D=1
M8 out_b 14 18 gnd! NMOS_VTL L=5e-08 W=2.7e-07 AD=3.105e-14 AS=3.78e-14 PD=7.7e-07 PS=8.2e-07 $X=6435 $Y=-935 $D=1
M9 4 A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=1.935e-14 PD=5.85e-07 PS=5.75e-07 $X=-705 $Y=3505 $D=0
M10 vdd! out 4 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=115 $Y=3505 $D=0
M11 6 !A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=900 $Y=3505 $D=0
M12 vdd! out_b 6 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=1720 $Y=3505 $D=0
M13 8 !B vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=2530 $Y=3505 $D=0
M14 vdd! out_b 8 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3305 $Y=3505 $D=0
M15 14 !C vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=4030 $Y=3505 $D=0
M16 vdd! out_b 14 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=4850 $Y=3505 $D=0
M17 out_b 6 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07 $X=5675 $Y=855 $D=0
M18 vdd! 8 out_b vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.52e-14 PD=6.4e-07 PS=6.4e-07 $X=6055 $Y=855 $D=0
M19 out_b 14 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=2.52e-14 PD=5.75e-07 PS=6.4e-07 $X=6435 $Y=855 $D=0
X20 4 gnd! vdd! out INV $T=6065 2910 0 0 $X=5615 $Y=2395
.ENDS
***************************************
.SUBCKT BE_Cell Yj+1_b Yj+1 Yj_b Yj Yj-1_b Yj-1 gnd! vdd! TWO TWO_b ONE_b ONE
** N=16 EP=12 IP=36 FDC=82
X0 TWO_b 11 TWO 9 gnd! vdd! 10 13 SP_OR_DR $T=36600 -5140 0 0 $X=36595 $Y=-5535
X1 Yj-1 ONE Yj-1_b ONE_b Yj gnd! vdd! Yj_b SP_XOR_DR $T=37070 -13205 0 0 $X=37070 $Y=-13600
X2 Yj+1_b Yj Yj-1 9 10 gnd! vdd! Yj+1 Yj_b Yj-1_b SP_AND3_DR $T=25560 -12380 0 0 $X=23610 $Y=-13600
X3 Yj+1 Yj_b Yj-1_b 11 13 gnd! vdd! Yj+1_b Yj Yj-1 SP_AND3_DR $T=25560 -5140 0 0 $X=23610 $Y=-6360
.ENDS
***************************************
.SUBCKT MULT_TOP_v1 vdd! gnd! VDD_PC GND_PC X15_b X15 X14_b X14 X13_b X13 X12_b X12 X11_b X11 X10_b X10 X9_b X9 Y15 Y15_b
+ X8_b X8 X7_b X7 X6_b X6 X5_b X5 X4_b X4 X3_b X3 X2_b X2 X1_b X1 X0_b X0 Y13_b Y13
+ Y11_b Y11 Y9_b Y9 Y7_b Y7 Y5_b Y5 Y3_b Y3 Y1_b Y1 Y14_b Y14 Y12_b Y12 Y10_b Y10 Y8_b Y8
+ Y6_b Y6 Y4_b Y4 Y2_b Y2 Y0_b Y0 OV S31 S30 S29 S28 S27 S26 S25 S24 S23 S22 S21
+ S20 S19 S18 S17 S16 S15 S14 S13 S12 S11 S10 S9 S8 S7 S6 S5 S4 S3 S2 S1
+ S0
** N=961 EP=101 IP=3257 FDC=29664
X726 vdd! 555 557 25 556 gnd! 558 26 559 560 gnd! gnd! SP_FA_DR $T=1370670 294245 0 0 $X=1374990 $Y=294745
X727 vdd! 567 569 27 568 gnd! 570 28 571 572 561 566 SP_FA_DR $T=1388630 294245 0 0 $X=1392950 $Y=294745
X728 vdd! 579 581 29 580 gnd! 582 30 583 584 573 578 SP_FA_DR $T=1406590 294245 0 0 $X=1410910 $Y=294745
X729 vdd! 591 593 31 592 gnd! 594 32 595 596 585 590 SP_FA_DR $T=1424550 294245 0 0 $X=1428870 $Y=294745
X730 vdd! 603 605 33 604 gnd! 606 34 607 608 597 602 SP_FA_DR $T=1442510 294245 0 0 $X=1446830 $Y=294745
X731 vdd! 615 617 35 616 gnd! 618 36 619 620 609 614 SP_FA_DR $T=1460470 294245 0 0 $X=1464790 $Y=294745
X732 vdd! 627 629 37 628 gnd! 630 38 631 633 621 626 SP_FA_DR $T=1478430 294245 0 0 $X=1482750 $Y=294745
X733 vdd! 641 643 39 642 gnd! 644 40 645 647 635 640 SP_FA_DR $T=1496390 294245 0 0 $X=1500710 $Y=294745
X734 vdd! 654 656 41 655 gnd! 657 42 658 660 648 653 SP_FA_DR $T=1514350 294245 0 0 $X=1518670 $Y=294745
X735 vdd! 668 670 43 669 gnd! 671 44 672 673 661 667 SP_FA_DR $T=1532310 294245 0 0 $X=1536630 $Y=294745
X736 vdd! 681 683 45 682 gnd! 684 46 685 686 674 680 SP_FA_DR $T=1550270 294245 0 0 $X=1554590 $Y=294745
X737 vdd! 694 696 47 695 gnd! 697 48 698 700 688 693 SP_FA_DR $T=1568230 294245 0 0 $X=1572550 $Y=294745
X738 vdd! 707 709 49 708 gnd! 710 50 712 713 701 706 SP_FA_DR $T=1586190 294245 0 0 $X=1590510 $Y=294745
X739 vdd! 721 723 52 722 gnd! 724 53 725 726 714 720 SP_FA_DR $T=1604150 294245 0 0 $X=1608470 $Y=294745
X740 vdd! 734 736 55 735 gnd! 737 56 738 739 728 733 SP_FA_DR $T=1622110 294245 0 0 $X=1626430 $Y=294745
X741 vdd! 747 749 57 748 gnd! 750 58 751 753 741 746 SP_FA_DR $T=1640070 294245 0 0 $X=1644390 $Y=294745
X742 vdd! 761 763 GND_PC 762 gnd! 764 VDD_PC 765 766 754 759 SP_FA_DR $T=1658030 294245 0 0 $X=1662350 $Y=294745
X743 vdd! 774 776 Y15 775 gnd! 777 Y15_b 778 779 767 773 SP_FA_DR $T=1675990 294245 0 0 $X=1680310 $Y=294745
X744 vdd! 787 789 GND_PC 788 gnd! 790 VDD_PC 791 793 781 786 SP_FA_DR $T=1693950 294245 0 0 $X=1698270 $Y=294745
X745 vdd! 800 802 GND_PC 801 gnd! 803 VDD_PC 805 806 794 799 SP_FA_DR $T=1711910 294245 0 0 $X=1716230 $Y=294745
X746 vdd! 814 816 GND_PC 815 gnd! 817 VDD_PC 818 819 807 813 SP_FA_DR $T=1729870 294245 0 0 $X=1734190 $Y=294745
X747 vdd! 827 829 GND_PC 828 gnd! 830 VDD_PC 831 832 821 826 SP_FA_DR $T=1747830 294245 0 0 $X=1752150 $Y=294745
X748 vdd! 840 842 GND_PC 841 gnd! 843 VDD_PC 844 846 834 839 SP_FA_DR $T=1765790 294245 0 0 $X=1770110 $Y=294745
X749 vdd! 853 855 GND_PC 854 gnd! 857 VDD_PC 858 859 847 852 SP_FA_DR $T=1783750 294245 0 0 $X=1788070 $Y=294745
X750 vdd! 867 869 GND_PC 868 gnd! 870 VDD_PC 871 872 860 866 SP_FA_DR $T=1801710 294245 0 0 $X=1806030 $Y=294745
X751 vdd! 880 882 GND_PC 881 gnd! 883 VDD_PC 884 886 874 879 SP_FA_DR $T=1819670 294245 0 0 $X=1823990 $Y=294745
X752 vdd! 893 895 GND_PC 894 gnd! 896 VDD_PC 897 899 887 892 SP_FA_DR $T=1837630 294245 0 0 $X=1841950 $Y=294745
X753 vdd! 907 909 GND_PC 908 gnd! 910 VDD_PC 911 912 900 906 SP_FA_DR $T=1855590 294245 0 0 $X=1859910 $Y=294745
X754 vdd! 920 922 GND_PC 921 gnd! 923 VDD_PC 924 925 913 919 SP_FA_DR $T=1873550 294245 0 0 $X=1877870 $Y=294745
X755 vdd! 933 935 GND_PC 934 gnd! 936 VDD_PC 937 939 927 928 SP_FA_DR $T=1891510 294245 0 0 $X=1895830 $Y=294745
X756 vdd! 946 948 GND_PC 947 gnd! 949 VDD_PC 950 954 940 941 SP_FA_DR $T=1909470 294245 0 0 $X=1913790 $Y=294745
X757 vdd! GND_PC 958 GND_PC VDD_PC gnd! 959 VDD_PC 960 961 952 953 SP_FA_DR $T=1927430 294245 0 0 $X=1931750 $Y=294745
X764 gnd! VDD_PC GND_PC gnd! 5 6 7 8 VDD_PC gnd! GND_PC vdd! X15_b X15 gnd! gnd! X14_b X14 25 26
+ X13_b X13 27 28 X12_b X12 29 30 X11_b X11 31 32 X10_b X10 33 34 X9_b X9 35 36
+ X8_b X8 37 38 39 40 41 42 43 44 45 46 47 48 49 50 52 53 55 56
+ X7_b 57 58 X7 X6_b X6 X5_b X5 X4_b X4 X3_b X3 X2_b X2 X1_b X1 X0_b X0
+ PPG_Blk_v1 $T=130430 503570 0 0 $X=164190 $Y=527855
X765 gnd! VDD_PC GND_PC 79 75 76 77 78 Y15_b 80 Y15 vdd! X15_b X15 81 82 X14_b X14 83 84
+ X13_b X13 85 86 X12_b X12 87 88 X11_b X11 89 90 X10_b X10 91 92 X9_b X9 93 94
+ X8_b X8 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112
+ X7_b 113 114 X7 X6_b X6 X5_b X5 X4_b X4 X3_b X3 X2_b X2 X1_b X1 X0_b X0
+ PPG_Blk_v1 $T=343220 503570 0 0 $X=376980 $Y=527855
X766 gnd! VDD_PC GND_PC 115 173 174 175 176 Y13_b 116 Y13 vdd! X15_b X15 117 118 X14_b X14 119 120
+ X13_b X13 121 122 X12_b X12 123 124 X11_b X11 125 126 X10_b X10 127 128 X9_b X9 129 130
+ X8_b X8 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148
+ X7_b 149 150 X7 X6_b X6 X5_b X5 X4_b X4 X3_b X3 X2_b X2 X1_b X1 X0_b X0
+ PPG_Blk_v1 $T=555945 503570 0 0 $X=589705 $Y=527855
X767 gnd! VDD_PC GND_PC 153 267 268 269 270 Y11_b 154 Y11 vdd! X15_b X15 181 182 X14_b X14 187 188
+ X13_b X13 195 196 X12_b X12 203 204 X11_b X11 211 212 X10_b X10 219 220 X9_b X9 227 228
+ X8_b X8 235 236 243 244 251 252 259 260 273 274 281 282 289 290 297 298 305 306
+ X7_b 313 314 X7 X6_b X6 X5_b X5 X4_b X4 X3_b X3 X2_b X2 X1_b X1 X0_b X0
+ PPG_Blk_v1 $T=768685 503570 0 0 $X=802445 $Y=527855
X768 gnd! VDD_PC GND_PC 151 349 350 351 352 Y9_b 152 Y9 vdd! X15_b X15 193 194 X14_b X14 201 202
+ X13_b X13 209 210 X12_b X12 217 218 X11_b X11 225 226 X10_b X10 233 234 X9_b X9 241 242
+ X8_b X8 249 250 257 258 271 272 279 280 287 288 295 296 303 304 311 312 319 320
+ X7_b 325 326 X7 X6_b X6 X5_b X5 X4_b X4 X3_b X3 X2_b X2 X1_b X1 X0_b X0
+ PPG_Blk_v1 $T=981385 503570 0 0 $X=1015145 $Y=527855
X769 gnd! VDD_PC GND_PC 373 369 370 371 372 Y7_b 374 Y7 vdd! X15_b X15 375 376 X14_b X14 377 378
+ X13_b X13 379 380 X12_b X12 381 382 X11_b X11 383 384 X10_b X10 385 386 X9_b X9 387 388
+ X8_b X8 389 390 391 392 393 394 395 396 397 398 399 400 401 402 403 404 405 406
+ X7_b 407 408 X7 X6_b X6 X5_b X5 X4_b X4 X3_b X3 X2_b X2 X1_b X1 X0_b X0
+ PPG_Blk_v1 $T=1194115 503570 0 0 $X=1227875 $Y=527855
X770 gnd! VDD_PC GND_PC 409 451 452 453 454 Y5_b 410 Y5 vdd! X15_b X15 411 412 X14_b X14 413 414
+ X13_b X13 415 416 X12_b X12 417 418 X11_b X11 419 420 X10_b X10 421 422 X9_b X9 423 424
+ X8_b X8 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ X7_b 443 444 X7 X6_b X6 X5_b X5 X4_b X4 X3_b X3 X2_b X2 X1_b X1 X0_b X0
+ PPG_Blk_v1 $T=1406840 503570 0 0 $X=1440600 $Y=527855
X771 gnd! VDD_PC GND_PC 447 465 466 467 468 Y3_b 448 Y3 vdd! X15_b X15 455 456 X14_b X14 457 458
+ X13_b X13 461 462 X12_b X12 471 472 X11_b X11 475 476 X10_b X10 479 480 X9_b X9 483 484
+ X8_b X8 487 488 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506
+ X7_b 507 508 X7 X6_b X6 X5_b X5 X4_b X4 X3_b X3 X2_b X2 X1_b X1 X0_b X0
+ PPG_Blk_v1 $T=1619580 503570 0 0 $X=1653340 $Y=527855
X772 gnd! VDD_PC GND_PC 445 523 524 525 526 Y1_b 446 Y1 vdd! X15_b X15 459 460 X14_b X14 469 470
+ X13_b X13 473 474 X12_b X12 477 478 X11_b X11 481 482 X10_b X10 485 486 X9_b X9 489 490
+ X8_b X8 509 510 511 512 513 514 515 516 517 518 519 520 527 528 529 530 531 532
+ X7_b 533 534 X7 X6_b X6 X5_b X5 X4_b X4 X3_b X3 X2_b X2 X1_b X1 X0_b X0
+ PPG_Blk_v1 $T=1832280 503570 0 0 $X=1866040 $Y=527855
X773 OV gnd! vdd! GND_PC S31 561 566 559 560 S30 573 578 571 572 S29 585 590 583 584 S28
+ 597 602 595 596 S27 609 614 607 608 S26 621 626 619 620 S25 635 640 631 633 S24
+ 648 653 645 647 S23 661 667 658 660 S22 674 680 672 673 S21 688 693 685 686 S20
+ 701 706 698 700 S19 714 720 712 713 S18 728 733 725 726 S17 741 746 738 739 S16
+ 754 759 751 753 S15 767 773 765 766 S14 781 786 778 779 S13 794 799 791 793 S12
+ 807 813 805 806 S11 821 826 818 819 S10 834 839 831 832 S9 847 852 844 846 S8
+ 860 866 858 859 S7 874 879 871 872 S6 887 892 884 886 S5 900 906 897 899 S4
+ 913 919 911 912 S3 927 928 924 925 S2 940 941 937 939 S1 952 953 950 954 VDD_PC
+ S0 GND_PC VDD_PC 960 961
+ PPA_v1 $T=1631420 36160 0 0 $X=1495060 $Y=63705
X774 gnd! vdd! 79 80 155 156 81 82 159 160 83 84 163 164 85 86 167 168 87 88
+ 177 178 89 90 183 184 91 92 189 190 93 94 197 198 95 96 205 206 97 98
+ 213 214 99 100 221 222 101 102 229 230 103 104 237 238 105 106 245 246 107 108
+ 253 254 109 110 261 262 111 112 275 276 113 114 283 284 GND_PC VDD_PC 291 292 Y13 Y13_b
+ 299 300 GND_PC VDD_PC 307 308 GND_PC VDD_PC 315 316 GND_PC VDD_PC 321 322 GND_PC VDD_PC 327 328 GND_PC VDD_PC
+ 331 332 GND_PC VDD_PC 335 336 GND_PC VDD_PC 339 340 GND_PC VDD_PC 343 344 GND_PC VDD_PC 353 354 GND_PC VDD_PC
+ 357 358 GND_PC VDD_PC 361 362 GND_PC VDD_PC 151 152 153 154 115 116 157 158 151 152 153 154
+ 115 116 161 162 151 152 153 154 115 116 165 166 151 152 153 154 117 118 169 170
+ 151 152 153 154 119 120 179 180 151 152 181 182 121 122 185 186 151 152 187 188
+ 123 124 191 192 193 194 195 196 125 126 199 200 201 202 203 204 127 128 207 208
+ 209 210 211 212 129 130 215 216 217 218 219 220 131 132 223 224 225 226 227 228
+ 133 134 231 232 233 234 235 236 135 136 239 240 241 242 243 244 137 138 247 248
+ 249 250 251 252 139 140 255 256 257 258 259 260 141 142 263 264 271 272 273 274
+ 143 144 277 278 279 280 281 282 145 146 285 286 287 288 289 290 147 148 293 294
+ 295 296 297 298 149 150 301 302 303 304 305 306 GND_PC VDD_PC 309 310 311 312 313 314
+ Y11 Y11_b 317 318 319 320 GND_PC VDD_PC GND_PC VDD_PC 323 324 325 326 Y9 Y9_b GND_PC VDD_PC 329 330
+ GND_PC VDD_PC GND_PC VDD_PC GND_PC VDD_PC 333 334 Y7 Y7_b GND_PC VDD_PC GND_PC VDD_PC 337 338 GND_PC VDD_PC GND_PC VDD_PC
+ GND_PC VDD_PC 341 342 GND_PC VDD_PC GND_PC VDD_PC GND_PC VDD_PC 345 346 GND_PC VDD_PC GND_PC VDD_PC GND_PC VDD_PC 355 356
+ GND_PC VDD_PC GND_PC VDD_PC GND_PC VDD_PC 359 360 GND_PC VDD_PC GND_PC VDD_PC GND_PC VDD_PC 363 364 GND_PC VDD_PC GND_PC VDD_PC
+ GND_PC VDD_PC 365 366
+ SP_42CSA_DR $T=623110 302395 0 0 $X=519290 $Y=429845
X775 gnd! vdd! 373 374 551 552 373 374 562 563 373 374 574 575 373 374 586 587 373 374
+ 598 599 373 374 610 611 373 374 622 623 373 374 636 637 373 374 649 650 375 376
+ 662 663 377 378 676 677 379 380 689 690 381 382 702 703 383 384 716 717 385 386
+ 729 730 387 388 742 743 389 390 755 756 391 392 769 770 393 394 782 783 395 396
+ 795 796 397 398 808 809 399 400 822 823 401 402 835 836 403 404 848 849 405 406
+ 862 863 407 408 875 876 GND_PC VDD_PC 888 889 Y5 Y5_b 901 902 GND_PC VDD_PC 915 916 GND_PC VDD_PC
+ 929 930 GND_PC VDD_PC 942 943 GND_PC VDD_PC 445 446 447 448 409 410 553 554 445 446 447 448
+ 409 410 564 565 445 446 447 448 409 410 576 577 445 446 447 448 409 410 588 589
+ 445 446 447 448 409 410 600 601 445 446 447 448 409 410 612 613 445 446 447 448
+ 409 410 624 625 445 446 447 448 409 410 638 639 445 446 447 448 409 410 651 652
+ 445 446 447 448 409 410 664 665 445 446 447 448 409 410 678 679 445 446 447 448
+ 411 412 691 692 445 446 447 448 413 414 704 705 445 446 455 456 415 416 718 719
+ 445 446 457 458 417 418 731 732 459 460 461 462 419 420 744 745 469 470 471 472
+ 421 422 757 758 473 474 475 476 423 424 771 772 477 478 479 480 425 426 784 785
+ 481 482 483 484 427 428 797 798 485 486 487 488 429 430 811 812 489 490 491 492
+ 431 432 824 825 509 510 493 494 433 434 837 838 511 512 495 496 435 436 850 851
+ 513 514 497 498 437 438 864 865 515 516 499 500 439 440 877 878 517 518 501 502
+ 441 442 890 891 519 520 503 504 443 444 903 904 527 528 505 506 GND_PC VDD_PC 917 918
+ 529 530 507 508 Y3 Y3_b 931 932 531 532 GND_PC VDD_PC GND_PC VDD_PC 944 945 533 534 Y1 Y1_b
+ GND_PC VDD_PC 955 956
+ SP_42CSA_DR $T=1474005 302395 0 0 $X=1370185 $Y=429845
X776 gnd! vdd! 157 158 555 556 161 162 567 568 165 166 579 580 169 170 591 592 179 180
+ 603 604 185 186 615 616 191 192 627 628 199 200 641 642 207 208 654 655 215 216
+ 668 669 223 224 681 682 231 232 694 695 239 240 707 708 247 248 721 722 255 256
+ 734 735 263 264 747 748 277 278 761 762 285 286 774 775 293 294 787 788 301 302
+ 800 801 309 310 814 815 317 318 827 828 323 324 840 841 329 330 853 854 333 334
+ 867 868 337 338 880 881 341 342 893 894 345 346 907 908 355 356 920 921 359 360
+ 933 934 363 364 946 947 365 366 551 552 553 554 155 156 557 558 562 563 564 565
+ 159 160 569 570 574 575 576 577 163 164 581 582 586 587 588 589 167 168 593 594
+ 598 599 600 601 177 178 605 606 610 611 612 613 183 184 617 618 622 623 624 625
+ 189 190 629 630 636 637 638 639 197 198 643 644 649 650 651 652 205 206 656 657
+ 662 663 664 665 213 214 670 671 676 677 678 679 221 222 683 684 689 690 691 692
+ 229 230 696 697 702 703 704 705 237 238 709 710 716 717 718 719 245 246 723 724
+ 729 730 731 732 253 254 736 737 742 743 744 745 261 262 749 750 755 756 757 758
+ 275 276 763 764 769 770 771 772 283 284 776 777 782 783 784 785 291 292 789 790
+ 795 796 797 798 299 300 802 803 808 809 811 812 307 308 816 817 822 823 824 825
+ 315 316 829 830 835 836 837 838 321 322 842 843 848 849 850 851 327 328 855 857
+ 862 863 864 865 331 332 869 870 875 876 877 878 335 336 882 883 888 889 890 891
+ 339 340 895 896 901 902 903 904 343 344 909 910 915 916 917 918 353 354 922 923
+ 929 930 931 932 357 358 935 936 942 943 944 945 361 362 948 949 GND_PC VDD_PC 955 956
+ GND_PC VDD_PC 958 959
+ SP_42CSA_DR $T=1476060 205055 0 0 $X=1372240 $Y=332505
X791 VDD_PC GND_PC VDD_PC GND_PC Y15_b Y15 gnd! vdd! 8 7 5 6 BE_Cell $T=107425 594020 0 0 $X=126365 $Y=580420
X792 Y15_b Y15 Y14_b Y14 Y13_b Y13 gnd! vdd! 78 77 75 76 BE_Cell $T=107425 608480 0 0 $X=126365 $Y=594880
X793 Y13_b Y13 Y12_b Y12 Y11_b Y11 gnd! vdd! 176 175 173 174 BE_Cell $T=107425 622940 0 0 $X=126365 $Y=609340
X794 Y11_b Y11 Y10_b Y10 Y9_b Y9 gnd! vdd! 270 269 267 268 BE_Cell $T=107425 637405 0 0 $X=126365 $Y=623805
X795 Y9_b Y9 Y8_b Y8 Y7_b Y7 gnd! vdd! 352 351 349 350 BE_Cell $T=107425 651870 0 0 $X=126365 $Y=638270
X796 Y7_b Y7 Y6_b Y6 Y5_b Y5 gnd! vdd! 372 371 369 370 BE_Cell $T=107425 666330 0 0 $X=126365 $Y=652730
X797 Y5_b Y5 Y4_b Y4 Y3_b Y3 gnd! vdd! 454 453 451 452 BE_Cell $T=107425 680790 0 0 $X=126365 $Y=667190
X798 Y3_b Y3 Y2_b Y2 Y1_b Y1 gnd! vdd! 468 467 465 466 BE_Cell $T=107425 695255 0 0 $X=126365 $Y=681655
X799 Y1_b Y1 Y0_b Y0 VDD_PC GND_PC gnd! vdd! 526 525 523 524 BE_Cell $T=107425 709720 0 0 $X=126365 $Y=696120
.ENDS
***************************************
