* SPICE NETLIST
***************************************

.SUBCKT INV in gnd! vdd! out
** N=4 EP=4 IP=0 FDC=2
M0 out in gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07 $X=210 $Y=-180 $D=1
M1 out in vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07 $X=210 $Y=800 $D=0
.ENDS
***************************************
.SUBCKT NAND2 A gnd! B OUT vdd!
** N=6 EP=5 IP=0 FDC=4
M0 6 A gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07 $X=210 $Y=-360 $D=1
M1 OUT B 6 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=2.52e-14 PD=5.75e-07 PS=6.4e-07 $X=590 $Y=-360 $D=1
M2 OUT A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07 $X=210 $Y=670 $D=0
M3 vdd! B OUT vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14 PD=5.7e-07 PS=6.4e-07 $X=590 $Y=670 $D=0
.ENDS
***************************************
.SUBCKT BLACK_CELL Pi-1 !Pi-1 Gi !Gi Pi !Pi !Gi-1 Gi-1 !G P G !P gnd! vdd!
** N=23 EP=14 IP=18 FDC=34
M0 22 Pi-1 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.025e-14 PD=6.4e-07 PS=5.85e-07 $X=690 $Y=10785 $D=1
M1 20 !Gi 9 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07 $X=1060 $Y=5725 $D=1
M2 10 Pi 22 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=2.52e-14 PD=6.65e-07 PS=6.4e-07 $X=1070 $Y=10785 $D=1
M3 20 !Gi-1 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07 $X=1930 $Y=5725 $D=1
M4 gnd! !Pi 20 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14 PD=5.7e-07 PS=6.4e-07 $X=2310 $Y=5725 $D=1
M5 13 !Pi gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=2320 $Y=10785 $D=1
M6 gnd! Gi 14 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3140 $Y=5725 $D=1
M7 23 Gi-1 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.88e-14 AS=2.025e-14 PD=6.8e-07 PS=5.85e-07 $X=3950 $Y=5725 $D=1
M8 21 !Pi-1 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3950 $Y=10785 $D=1
M9 17 Pi 23 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.385e-14 AS=2.88e-14 PD=6.25e-07 PS=6.8e-07 $X=4370 $Y=5725 $D=1
M10 9 !Gi vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=690 $Y=9120 $D=0
M11 10 Pi vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=690 $Y=14180 $D=0
M12 vdd! !G 9 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=1510 $Y=9120 $D=0
M13 vdd! P 10 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=1510 $Y=14180 $D=0
M14 14 Gi vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=2320 $Y=9120 $D=0
M15 13 !Pi vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=2320 $Y=14180 $D=0
M16 vdd! G 14 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3140 $Y=9120 $D=0
M17 vdd! !P 13 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3140 $Y=14180 $D=0
M18 17 Pi vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=3950 $Y=9120 $D=0
M19 21 !Pi-1 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=3950 $Y=14180 $D=0
M20 vdd! G 17 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=4770 $Y=9120 $D=0
M21 vdd! !P 21 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=4770 $Y=14180 $D=0
X22 10 gnd! vdd! P INV $T=6080 13585 0 0 $X=5630 $Y=13070
X23 9 gnd! vdd! !G INV $T=6620 5735 0 0 $X=6170 $Y=5220
X24 14 gnd! 17 G vdd! NAND2 $T=6200 8655 0 0 $X=5750 $Y=8010
X25 21 gnd! 13 !P vdd! NAND2 $T=6270 10925 0 0 $X=5820 $Y=10280
.ENDS
***************************************
