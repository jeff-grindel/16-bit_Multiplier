* SPICE NETLIST
***************************************

.SUBCKT NAND2 A gnd! B OUT vdd!
** N=6 EP=5 IP=0 FDC=4
M0 6 A gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07 $X=210 $Y=-360 $D=1
M1 OUT B 6 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=2.52e-14 PD=5.75e-07 PS=6.4e-07 $X=590 $Y=-360 $D=1
M2 OUT A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07 $X=210 $Y=670 $D=0
M3 vdd! B OUT vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14 PD=5.7e-07 PS=6.4e-07 $X=590 $Y=670 $D=0
.ENDS
***************************************
.SUBCKT SP_XOR P !A B !B A gnd! vdd!
** N=11 EP=7 IP=5 FDC=12
M0 10 !B gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.025e-14 PD=6.4e-07 PS=5.85e-07 $X=675 $Y=110 $D=1
M1 1 A 10 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=2.52e-14 PD=6.65e-07 PS=6.4e-07 $X=1055 $Y=110 $D=1
M2 11 !A 3 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.745e-14 PD=6.4e-07 PS=6.65e-07 $X=2745 $Y=110 $D=1
M3 gnd! B 11 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.52e-14 PD=5.85e-07 PS=6.4e-07 $X=3125 $Y=110 $D=1
M4 1 A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=675 $Y=2740 $D=0
M5 vdd! P 1 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=1495 $Y=2740 $D=0
M6 3 P vdd! vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=2305 $Y=2740 $D=0
M7 vdd! !A 3 vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=3125 $Y=2740 $D=0
X8 1 gnd! 3 P vdd! NAND2 $T=4925 470 0 0 $X=4475 $Y=-175
.ENDS
***************************************
.SUBCKT INV in gnd! vdd! out
** N=4 EP=4 IP=0 FDC=2
M0 out in gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07 $X=210 $Y=-180 $D=1
M1 out in vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07 $X=210 $Y=800 $D=0
.ENDS
***************************************
.SUBCKT SP_AND_DR out !A out_b !B gnd! vdd! B A
** N=12 EP=8 IP=9 FDC=16
M0 12 B gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.025e-14 PD=6.4e-07 PS=5.85e-07 $X=675 $Y=110 $D=1
M1 1 A 12 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=2.52e-14 PD=6.65e-07 PS=6.4e-07 $X=1055 $Y=110 $D=1
M2 4 !A gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=2305 $Y=110 $D=1
M3 11 !B gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3935 $Y=110 $D=1
M4 1 A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=675 $Y=3505 $D=0
M5 vdd! out 1 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=1495 $Y=3505 $D=0
M6 4 !A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=2305 $Y=3505 $D=0
M7 vdd! out_b 4 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3125 $Y=3505 $D=0
M8 11 !B vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=3935 $Y=3505 $D=0
M9 vdd! out_b 11 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=4755 $Y=3505 $D=0
X10 11 gnd! 4 out_b vdd! NAND2 $T=6255 250 0 0 $X=5805 $Y=-395
X11 1 gnd! vdd! out INV $T=6065 2910 0 0 $X=5615 $Y=2395
.ENDS
***************************************
.SUBCKT PG_Blk !A A B !B P !P gnd! vdd! !G G
** N=16 EP=10 IP=18 FDC=38
M0 5 !B gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.025e-14 PD=6.4e-07 PS=5.85e-07 $X=2175 $Y=8750 $D=1
M1 6 A 5 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=2.52e-14 PD=6.65e-07 PS=6.4e-07 $X=2555 $Y=8750 $D=1
M2 8 !A 5 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=5.445e-14 PD=6.65e-07 PS=9.65e-07 $X=4185 $Y=8750 $D=1
M3 10 B gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.025e-14 PD=6.4e-07 PS=5.85e-07 $X=5455 $Y=8750 $D=1
M4 11 !A 10 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=2.52e-14 PD=6.65e-07 PS=6.4e-07 $X=5835 $Y=8750 $D=1
M5 14 A 10 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=5.445e-14 PD=6.65e-07 PS=9.65e-07 $X=7465 $Y=8750 $D=1
M6 6 A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=2175 $Y=12145 $D=0
M7 vdd! P 6 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=2995 $Y=12145 $D=0
M8 8 !A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=3805 $Y=12145 $D=0
M9 vdd! !P 8 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=4625 $Y=12145 $D=0
M10 11 !A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=5455 $Y=12145 $D=0
M11 vdd! P 11 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=6275 $Y=12145 $D=0
M12 14 A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=7085 $Y=12145 $D=0
M13 vdd! !P 14 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=7905 $Y=12145 $D=0
X14 14 gnd! 8 !P vdd! NAND2 $T=9320 8890 0 0 $X=8870 $Y=8245
X15 6 gnd! 11 P vdd! NAND2 $T=9320 11680 0 0 $X=8870 $Y=11035
X16 G !A !G !B gnd! vdd! B A SP_AND_DR $T=1500 3355 0 0 $X=1495 $Y=2960
.ENDS
***************************************
.SUBCKT GREY_CELL !Gi-1 Gi-1 !Gi Gi !Pi Pi !G G gnd! vdd!
** N=15 EP=10 IP=9 FDC=18
M0 14 !Gi 7 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07 $X=1045 $Y=110 $D=1
M1 14 !Gi-1 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07 $X=1915 $Y=110 $D=1
M2 gnd! !Pi 14 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14 PD=5.7e-07 PS=6.4e-07 $X=2295 $Y=110 $D=1
M3 gnd! Gi 9 gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3125 $Y=110 $D=1
M4 15 Gi-1 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.88e-14 AS=2.025e-14 PD=6.8e-07 PS=5.85e-07 $X=3935 $Y=110 $D=1
M5 11 Pi 15 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.385e-14 AS=2.88e-14 PD=6.25e-07 PS=6.8e-07 $X=4355 $Y=110 $D=1
M6 7 !Gi vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=675 $Y=3505 $D=0
M7 vdd! !G 7 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=1495 $Y=3505 $D=0
M8 9 Gi vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=2305 $Y=3505 $D=0
M9 vdd! G 9 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3125 $Y=3505 $D=0
M10 11 Pi vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=3935 $Y=3505 $D=0
M11 vdd! G 11 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=4755 $Y=3505 $D=0
X12 9 gnd! 11 G vdd! NAND2 $T=6185 3040 0 0 $X=5735 $Y=2395
X13 7 gnd! vdd! !G INV $T=6605 120 0 0 $X=6155 $Y=-395
.ENDS
***************************************
.SUBCKT BLACK_CELL Pi-1 !Pi-1 Gi !Gi Pi !Pi !Gi-1 gnd! vdd! Gi-1 !G G !P P
** N=14 EP=14 IP=18 FDC=34
X0 P !Pi !P !Pi-1 gnd! vdd! Pi-1 Pi SP_AND_DR $T=15 10675 0 0 $X=10 $Y=10280
X1 !Gi-1 Gi-1 !Gi Gi !Pi Pi !G G gnd! vdd! GREY_CELL $T=15 5615 0 0 $X=0 $Y=5220
.ENDS
***************************************
.SUBCKT PPA4 vdd! gnd! S3 A3 A3_b B3 B3_b S2 A2 A2_b B2 B2_b S1 A1 A1_b B1 B1_b S0 A0 A0_b
+ B0 B0_b
** N=51 EP=22 IP=126 FDC=322
X0 S3 3 4 5 2 gnd! vdd! SP_XOR $T=264770 150340 1 270 $X=261165 $Y=143940
X1 S2 8 10 12 7 gnd! vdd! SP_XOR $T=278820 150340 1 270 $X=275215 $Y=143940
X2 S1 14 16 18 13 gnd! vdd! SP_XOR $T=295545 150340 1 270 $X=291940 $Y=143940
X3 S0 19 gnd! vdd! 46 gnd! vdd! SP_XOR $T=309595 150340 1 270 $X=305990 $Y=143940
X4 A3_b A3 B3 B3_b 2 3 gnd! vdd! 31 25 PG_Blk $T=277700 210235 1 270 $X=264690 $Y=198830
X5 A2_b A2 B2 B2_b 7 8 gnd! vdd! 11 9 PG_Blk $T=291750 210235 1 270 $X=278740 $Y=198830
X6 A1_b A1 B1 B1_b 13 14 gnd! vdd! 17 15 PG_Blk $T=305800 210235 1 270 $X=292790 $Y=198830
X7 A0_b A0 B0 B0_b 46 19 gnd! vdd! 18 16 PG_Blk $T=319850 210235 1 270 $X=306840 $Y=198830
X8 12 10 30 29 27 26 gnd! gnd! gnd! vdd! GREY_CELL $T=274235 169410 1 270 $X=269865 $Y=161075
X9 18 16 40 39 37 36 5 4 gnd! vdd! GREY_CELL $T=288285 169410 1 270 $X=283915 $Y=161075
X10 18 16 17 15 14 13 12 10 gnd! vdd! GREY_CELL $T=302445 192410 1 270 $X=298075 $Y=184075
X11 7 8 25 31 2 3 11 gnd! vdd! 9 30 29 27 26 BLACK_CELL $T=279850 189975 1 270 $X=264805 $Y=181375
X12 13 14 9 11 7 8 17 gnd! vdd! 15 40 39 37 36 BLACK_CELL $T=293900 189975 1 270 $X=278855 $Y=181375
.ENDS
***************************************
