* SPICE NETLIST
***************************************

.SUBCKT INV in gnd! vdd! out
** N=4 EP=4 IP=0 FDC=2
M0 out in gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07 $X=210 $Y=-180 $D=1
M1 out in vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07 $X=210 $Y=800 $D=0
.ENDS
***************************************
.SUBCKT NAND2 A gnd! B OUT vdd!
** N=6 EP=5 IP=0 FDC=4
M0 6 A gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07 $X=210 $Y=-360 $D=1
M1 OUT B 6 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=1.935e-14 AS=2.52e-14 PD=5.75e-07 PS=6.4e-07 $X=590 $Y=-360 $D=1
M2 OUT A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07 $X=210 $Y=670 $D=0
M3 vdd! B OUT vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14 PD=5.7e-07 PS=6.4e-07 $X=590 $Y=670 $D=0
.ENDS
***************************************
.SUBCKT SP_AND_DR out !A out_b !B gnd! vdd! B A
** N=12 EP=8 IP=9 FDC=16
M0 12 B gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.025e-14 PD=6.4e-07 PS=5.85e-07 $X=675 $Y=110 $D=1
M1 1 A 12 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=2.52e-14 PD=6.65e-07 PS=6.4e-07 $X=1055 $Y=110 $D=1
M2 4 !A gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=2305 $Y=110 $D=1
M3 11 !B gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3935 $Y=110 $D=1
M4 1 A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=675 $Y=3505 $D=0
M5 vdd! out 1 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=1495 $Y=3505 $D=0
M6 4 !A vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=2305 $Y=3505 $D=0
M7 vdd! out_b 4 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=3125 $Y=3505 $D=0
M8 11 !B vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=3935 $Y=3505 $D=0
M9 vdd! out_b 11 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=4755 $Y=3505 $D=0
X10 1 gnd! vdd! out INV $T=6065 2910 0 0 $X=5615 $Y=2395
X11 11 gnd! 4 out_b vdd! NAND2 $T=6255 250 0 0 $X=5805 $Y=-395
.ENDS
***************************************
.SUBCKT PPG_Cell POS_b POS TWO_b TWO Xj-1 Xj-1_b ONE_b Xj_b Xj vdd! gnd! PPG PPG_b ONE
** N=30 EP=14 IP=35 FDC=70
M0 30 27 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.025e-14 PD=6.4e-07 PS=5.85e-07 $X=16655 $Y=16685 $D=1
M1 14 12 30 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=2.52e-14 PD=6.65e-07 PS=6.4e-07 $X=17035 $Y=16685 $D=1
M2 16 11 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=18285 $Y=16685 $D=1
M3 28 13 gnd! gnd! NMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=19915 $Y=16685 $D=1
M4 19 15 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.025e-14 PD=6.4e-07 PS=5.85e-07 $X=26270 $Y=16685 $D=1
M5 20 POS 19 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=2.52e-14 PD=6.65e-07 PS=6.4e-07 $X=26650 $Y=16685 $D=1
M6 22 POS_b 19 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=5.445e-14 PD=6.65e-07 PS=9.65e-07 $X=28280 $Y=16685 $D=1
M7 24 17 gnd! gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=2.025e-14 PD=6.4e-07 PS=5.85e-07 $X=29550 $Y=16685 $D=1
M8 25 POS_b 24 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=2.52e-14 PD=6.65e-07 PS=6.4e-07 $X=29930 $Y=16685 $D=1
M9 29 POS 24 gnd! NMOS_VTL L=5e-08 W=1.8e-07 AD=2.745e-14 AS=5.445e-14 PD=6.65e-07 PS=9.65e-07 $X=31560 $Y=16685 $D=1
M10 14 12 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=16655 $Y=20080 $D=0
M11 vdd! 15 14 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=17475 $Y=20080 $D=0
M12 16 11 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=18285 $Y=20080 $D=0
M13 vdd! 17 16 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=19105 $Y=20080 $D=0
M14 28 13 vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=19915 $Y=20080 $D=0
M15 vdd! 17 28 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=20735 $Y=20080 $D=0
M16 20 POS vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=26270 $Y=20080 $D=0
M17 vdd! PPG 20 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=27090 $Y=20080 $D=0
M18 22 POS_b vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=27900 $Y=20080 $D=0
M19 vdd! PPG_b 22 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=28720 $Y=20080 $D=0
M20 25 POS_b vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=29550 $Y=20080 $D=0
M21 vdd! PPG 25 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=30370 $Y=20080 $D=0
M22 29 POS vdd! vdd! PMOS_VTL L=5e-08 W=1.8e-07 AD=2.025e-14 AS=2.025e-14 PD=5.85e-07 PS=5.85e-07 $X=31180 $Y=20080 $D=0
M23 vdd! PPG_b 29 vdd! PMOS_VTL L=5e-08 W=9e-08 AD=1.0125e-14 AS=1.0125e-14 PD=4.05e-07 PS=4.05e-07 $X=32000 $Y=20080 $D=0
X24 14 gnd! vdd! 15 INV $T=22045 19485 0 0 $X=21595 $Y=18970
X25 28 gnd! 16 17 vdd! NAND2 $T=22235 16825 0 0 $X=21785 $Y=16180
X26 29 gnd! 22 PPG_b vdd! NAND2 $T=33415 16825 0 0 $X=32965 $Y=16180
X27 20 gnd! 25 PPG vdd! NAND2 $T=33415 19615 0 0 $X=32965 $Y=18970
X28 11 TWO_b 12 Xj-1_b gnd! vdd! Xj-1 TWO SP_AND_DR $T=6270 10385 0 0 $X=6265 $Y=9990
X29 13 ONE_b 27 Xj_b gnd! vdd! Xj ONE SP_AND_DR $T=6270 16575 0 0 $X=6265 $Y=16180
.ENDS
***************************************
